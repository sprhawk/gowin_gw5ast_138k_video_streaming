--
--Written by GowinSynthesis
--Tool Version "V1.9.11.02"
--Sun Sep 14 11:26:49 2025

--Source file index table:
--file0 "\/home/hongbo/.local/Gowin_V1.9.11.02_SP1_linux/IDE/ipcore/TSE_MAC/data/eth_mac_top.v"
--file1 "\/home/hongbo/.local/Gowin_V1.9.11.02_SP1_linux/IDE/ipcore/TSE_MAC/data/eth_mac.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
s7S00I1BZx/SbROGAXvg67ZWORLGvVEhr3NKsaVysWvXWAUzg/uFuZX/3Jl8gZuJzi5rPKvGZUmr
u2j/WzapALKSvyVIru2rU04KBteb7gYUkP0KeoxfA5HQS9WrTryqU84w6FZkCf1HOe1tbB39DV3d
OSEbv3UNX6b66h6vkK8TqMEwoqIhxhb7g9qx+KMSM8X/iKyPZZ+uPtKqxsnxr7knNMDS95sWFr/h
HYmbVZ6zBqHTHuRhIFi70bdoKmshoZAsuKtPEr4wUEWa3oUxzP/lLZVH6S2mXA6j5Vuab44brpdN
raxdu6VJ0FvZhVbBqvfHAkEC5mXmJyx4SXCNEw==

`protect encoding=(enctype="base64", line_length=76, bytes=453376)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
qDZ6ehWwS3TOSA4jN/ppiNYLJUU7X9voIAZaFfLHNwWy7Cyug8azNRga1YQKp+h8nRTinupvDNKS
G2kqVzwmGNZlZ2ANmFMp5QTRZ6q0z2Rar8bFGpuscPdr6pDDHVDySGfN6FaGKFhWOpXcwRsbZS+S
fWMEilQqa26HVBCKbUvkLtObuhQefNUh1NkzMh0ijL/qqJrN1bf4hw45Eff2AqO5IxLVRvys7zAU
Q4hSgBgZPeHPHpzcPTU085PnNp/V0CLpVEeR8vUE68tvJSYPVc3+RbERaVIhwIdrTpnSmeSmBrsu
ah3TJYjDDNo+iPbDDX/iWCY19TEtlxb6SaZL2uaNXrbVoYD+SZIQsja3hP648T0OgZMTyEFwzZW8
k4BYsSt1wjY9rQ5f9yD4E1GwcdEpBnXQ0ufOcgtEla2I9J8aKmcVfA0JSSkVOnu95+xiUTNxfTIK
vIeJeHNGhQj51UVsTSC5bFXROEz0wTlOLZN2U2o1UD/20mvsTdczXrnq3MPpq8bumDbcThcxNIdC
CcjeHwkqzqn+62wrI3GWOYY6oeUKRBzquBC5Z6PS8np0kWFGtd2yCEA+MNISnO3mDnD4HI3swn8A
iAhVbinGMw3AU0gxWnHbPhPsRQM8Otcb3pBTDcowUVZtWo5JRHRAjaxidj8OhWU4rVfqKteimVyh
UB0jUVRaeE4w7eoPefcoY3oe92EW58RCr6LVWbf9JXFGbc9O3rBZz3t+eEFf/uRuv3s4Pg1j5vEs
cAg8UVWY5ubKuLPIEf7Oueb4W/vbFGHNmaLMMtRKfhRegeuifEgw2/Nnu6b23CI+UtTu6xvnvvZO
WPyhRFYMkoFu6Q5229Rhmda4xzYK+ALxmddqU9p+qKTLliCmdYiCwcUeFnyJNhWBiEZpJd8lPlzj
TUksK9ciusRQEi+Q+EoJEJFb1Z44Zf89K+Ba3X7wk0rcfVbp8KzgXKdYHr+rYIjK7DUop9rW3zlT
Ed4gTJqjBfagwKY+pLFzRzu9IvQdEYRijauhvIhVYSYTqHDDC/FKEbIXcTnNOqhjHhWfsBOkpyFv
Gk1LTSQajcvFhLE2VEpqa5/ANdCwe9zDhmuI07X2NADszHkB18sl2WPpa1EjHFNACrdWaUnT1Non
+Td1oXJ9frgJMIjUvaujrzrhF1IKogIDAh0DrIn66b3FGVCSciOakEH5UsfG2x52XaR1glNYFj6o
I2tRNind8LQl+16dp/xFyG83kvbV4tOrkJbJGOAGa92XFrHCM2s+p//G2PN9EezF/vtPUns7GKrs
Bg5gRpi4fyr7weHAFXYhOn0toIuXMnQqjb36NYZVF8EAAlQ21sHYr+fXLF+Lt7V473PYY5fQ+FTH
RTyd7PrwzJw5fXlaSa/bE7FrMPiIofP3HdpI8MYZGSP/J5KXa2ytqKF6zKpkxmnLj8yRQrGq1diE
bu2LkFyGddqS48VjZSTWpgbKVaD3ldNu2CYgn1yQ5SwdC6/AtZLwul0AKH+HKAzdAPZgPLpYnbSi
gwtBqL1JXzLDhLQ5kJKHRr4KgXL8IQtyLXn+22seErHNI6Yg6rVPTFDPA0GyKjeB78wEGmjWljeS
g61Xe2kpnCrxfgJaU0x+WxY7PS8K8IxSd/4GydGs9QJuuA1WAdM3PbIsKOJXNAoaDVtA4bjXD+Y4
m8siOlA+a0I6Tmc7dA2LiVK+sZjNHxrgK6GQOcZc7WD16m9ACfJcelkltQVniSV62yOvHV7azliy
jok34y3CFhZoAFtwNe8hSso3u8vdxR1eT1NneiQvgb5h9mKK58UsjMLYVJlZJj2jv/PMw/x1XAT3
WNNI2TUKbJIjr56vOespGPSKYetJHgaNZG9p/5Yn/ePs1XD1C3dgrYT9uCaX23WtHHKjeZHNOxh1
8fT6dhlJukmtZ4bDYqIbiHXFpK091S6hBn9w1KobrD02ZWA8TwW2z6STW/gM3cAWhk8TJA8JxeHe
cQC9VoXku9H2MD6nOMcNcIDLIRB1MrbHVZk+UnBI9AYpfKz7zrfWUVsc1hz9FhHxzSC4zItsGxZY
avDLhqtguDTgDknk2YFOqHmIYqep0I4RMbepXvVnltwCsCC8CLxSFLJ3GJ4HAVYvyx8r3Sh1If/z
bHCB6+X04lxv3oG5hFJHwtyIVuSwg+lXwz2xNUsUl2Ppc6HSzWb9ghq9Z42HyiZghl1Xkl4UrKk9
B3zKOTuFl4SXAYB63pAz0Mwucw6BblPWumOWoZ6OHC4BOAoaownGKqbmW2U9+i0R5vP9fpGn7ETV
tWEDNXEZuYfcocoHorrs75ftgAtoj5EysHJgZo0rwZwC9qrUeGi6yYocfsqk+EguXuivuDn5iIz2
zQ0/ZXzcAhmP4oy1k4Il6c4ojqPdHw8fFWgJ+cd4DFDYu+5mDFuBgh5PKLxKCU+4zbKLGqLbIdCV
Grhz0wfXtKzPOmHSIe0qe+NLBPoeesJJYQr3sn08zMiHvlJkU4yKTAMInOp+nqEQKuWO28H7CxAk
6jRQp1MlnXLkYHLgmuEQgu57EtNB4dzmpnMjs/2kv2gDml9LbzPn2IPx6hLlflKwmEDs0mdGLi9n
nzPZPQglSe/CC2WhEYY2n5ODts1BUg06P36IOlLvA+nJBBtHD8KqxkmDCEYjkEW1SgJMWx2VwefR
RW3Kv1oQapqJL8dB/neNTa/KplWF8PE8yfOLxewxEVBkTC6iSHFG/dWBxxKi47AFuCggu+bO0m5e
GTFH+gloRtHfJzkLPBcMHLwipCf7DHEZ9kQkHNxknXCSWt4Np/bvG/H1gh5vocTxParOA6dAn9EP
zfYoWrFVvi/X7+LLfBsJT/LXYvpteIL+o2vAID7lvJdaa/DJPxNADkxsA31jDZZJqZV1HcoocC5W
3v64B3BhCVUGZHQ3h/ixc5nnlX0xw8TClTOWuf5Uymvxhppq6YENDIMMqbbhgbosbmj2NpQfz5rp
Qn+N3FARPvi1RRKtkRHd4KfF5b1H+rP40noNBmwfWeH/ceDam9up7yksfHrlBJQA5qNTvSbREwcp
vBpraGp464MtLK+7Vz4Vvl3mXbW5fsTccHcbGCRRQtN/8kEf8qB8v2X2SOdiaOlsdrheu2WJKkaj
pD3WGXw9aInwykvecVuPNB8IkNP/nCPqZkha5xVFR7r1BV36YxXwiB12hid8r81JCJpLUpPweDt7
aL7MX7pysW4WKrACW/2m8+yoxSVjnmmx9RBeCA4kUGdbsYtP24P2sBtTTB2qZeo1RQE/GIasXf7U
YYsWwN/QJFtIJkRO8SmdAqeIXXEpDBI/3fTlaZ4gUUCtmg9hAkhb7wzuOxj4d2UkzmeSLJ4Vimmq
hu8cydcbn4hsGELtTrYonSXvCFqd+Ytl5HiIHmqYmpK8/GJbVZNlonMhc5wAB1UiWCMyZH8epPyS
2F8eYHKsqsH1F66echYk68bT/WVQ2iVO94FZi7bjtqZU9XxAzbcQGek2rPHhjvj/qzV9ZphsKp5P
bBo0QjUVHtzil9EH0h2AKooOZaMxUyAGijkfivpkR/FTntxoCdrtu90i5XnBG1K2Ff6ZTsrwH7ac
UCbdUbYTv4wppjDH+EdtxS0NeM5IhupEWgXLfFL9VZxOfpTY8fT2c7lUYKB3Fc5UjSIxXf6T64aV
UmVDuBaaUDIoEAExYj8SH0N6lSKXx9tnMH40x5+vGnprFKbKaL0yIiEVDAC627a2N34S2xxwiEiJ
F6oxFZC3jQQWXYZlc+4Gsd2fgNLciDwCPH2i+qhuAXbvHdGOMH2JSWaeImRjOj4VP31oO5IuzGum
f6+EylG5EVXcnksAi7yiDJoJzb30hbit9veWimoQUwLpmUlTSwdjhABNMqIdTKwReIz9rh+Y/MmD
SLD1R16idSiHc9YWgqhuSwXtukPJJoFES0RMtR2QlBucCqyLnA/04rMY+b4M7LvzA9ZLxFJ2QVMg
AzA2DWXQlaHzXFK5fbxdkCxN9P2EhK8nlAzzjSHLNNL6vCZWurguSMOPLEyrbFM6C6I9tbWv7o0A
D+eh9RyYtILhSLUm232QQ0oihtpcSlnACurJtYcwm4aoXXj8/Oou3jDL/9MUNwFeKoaCMjtARSuH
BDv8TEXulJZdOzt9bp9wyEcE3Ec315lxBsQKNFic9dWy3W3JuC1SfEs8rNwlnndBBNi3jF1a9PJx
LiIDwXeHx1FJwkskhiOTJLxA6KqtZDOwimjUy6+AQSyUzwCe1W7FOT1R4EF92vqM5XbpTOM1TX2x
c1lsay2u2XvPVIiRBamI70MsYGrtVu/yQz/TaThYFIWJQ2/XTcSXi25a5ZXidj16+P/8AAcTGukz
tYp7iHIjxYXLWGqgIrFci5wTKnQJO+CvyZ1AtBGYWgQwlMGDwo0s9RB8rjefpqEhGR2/RgwWdJt8
Iin0en0Mrzs70PAzdUoSZQsaVrXPkfMQUpRHHlfsmjEhf3l1KddA0VnCWY9N5TbmcZDEhsLUqkfh
T3zIVl9bodBeOwow6hS06vS7jL5VdRpj0qd7oTJ8BSouNA9Z6i+T+ZtHcuNGCuR3eE0lhRnlEwPu
WiYaaa2j7aeIe231sY0MN1FLtblJZhLy7FxfUEWOJtQjb41lQCkekfoXzTkkymihZ4oY+Bc8TWzN
fJoGGCbeLNp+B254H35G3k+wUZQO60gF9Za802Wmj7bUTuKdJpSgeJfUFFcN2p1IAjLHNhM/1jQ4
6PwIinHv/Rw0JKY5O3Zb5n+5GHjgZs8Jm20QIcYgWTbQHKUHzhOu5J5POyTU1KnhJeixKMP4myzb
6SJs2IOd6f4uTRLttGppIlyNgNmIGTU4j/P9OMS0tHYVUgT2Hk2Od6DQ7Z2nyrePgvdklXz+BvOX
yW9N4NBBpTU6NM7Ie9TPP4cYB915l6SCB/FA/EoH1/yCM6xH0a25XZxf9zvRsfPu3/UZKTZeQfhA
Z0PtZ430vzHHkRgLBnctaeGLj71/1zHTXxRBaZtUnpsqOotBzZ+X9tKNB0zoZES+NubDRMUhq1JD
5X9uPVI8cOhZcLSUAzeMhtbmLPFmoZ7qyW1S3WfmZr7TWWwEbMspv2e5ddU47tAip2JTlgkNFE/T
sH46G2ifq9fFQc5d5N3A0pj0jNYzlskXUwL0HRucrzKGiWhNIeIjFClWQCgMjjyO4JYm52d4+x0b
gVrufmy4Vcpzge0z7h5Y/s02xrsHPcKKWk3bfoedekWLWt/70NIsAh4pvBSsEyQ8SdXQFuHlf/Qe
EL9dd25yaHtDsX0Kf3P8M0jQLHwndc7+DC5GVQe2Npf2uJ1zpKrXeK79k2LxY83xduqE1+FNkNoM
lTi8WA00XJI1xyH+pw8AJ/oVeavyI5hPP8wYtwxyvaKIH6kRP2cFVNLQH6SvB34x6Z6xNA6SCiFe
hXxILLBYIxQ1xtpAXhkotDhL+OEzlyDmS8sPkC13zaK3pbfGP2++soCBRPTbO7CQykWfDgGOPe5A
448O5g7hn8A4lhW5MCvNphkJRcLxt5ylkQDBhsrAxbGNAR7an9hkNQLRonhX7VXjGTqNEyWpXcyW
PkabqP/kV+3i5RXV1eO40ZFMK0pu69qEy0FyHJek4VO5jxw0hyTa6X9zLmWqEc7M1EkrhFetbzVg
99viQIL0aki5qIViaR9G/PgCz3+aELDhrqJAEjbaHWwRvMbE6wSzYfSoBt/SQ93eV+0umj4dpc4O
Krjpglu159xx/4KB1dYgIzNp9cZ3o/jv+sLhWREa2aWRhCFewjTUTZJj6h+4k9bh0mgQlzwbg7qX
v//XNViz+3wdst4isn6qdHWezCpWFUdwWRQoioqjtvRJ4qwitJEP9C8CiBJVuMyD0+5CsespAyGQ
eem/pzmKo+WSd5vY3rUZMvNEMJgJFlnZxy7YCxGAM1NMn64QCYiuAhxVnzs5fEmg0Wi0L/KD22++
q57I6bwr2IrUvwmz4K5T54XNkLCBXPWbTdxL05TlMNNHJETaBlo14ohbRkKif2r8pg/W6Qw+E7ZM
YfMzuuNXHLMhV623QpTzzA0oZ+wbbwg+HouTSjFC+Yyqej7Sbl3WeTEq/c7z2anpWtihO4r9FIRI
0/hjrcFQI8VBUX71vMD1g8bREi8eDOXZ41S9PkDol7biTz4jRwJtNs0D8yRyG7e2B/XQpxJc3xv9
sxm8xDfpwrAiDCMkSzS5qPo87DvEl6BxVyaGrZn+fCQUBEGLKsAKAQhHF+xZtS2wOvN2tiZ0YmRU
ZjxNmE+BXbiIy795JP4b3HNtol2i5xIVDZyDsRwaOA/ELBCjLX4NP6MeOkVzpSpVXQi1OI1vKWJN
GXa1KOiyNGgOFTcy9tcYpwPe+WxCckl1RfVmTsCcPSQ+mfDderSzWbmXsOHYi+swrNMfxiL1tejU
WyK4oG+cwjTnw9mDDX6AlBEXBdPPbP7xwBcebSGxz3YucRpQRK8jssMiBN66nu/ncgOuQdbeiIOE
uCRWmDwM8izZM+LUt7gu86fZodBxR+4VU+PVfgHBpODdJWHxx6HbQ7lN62QfowoWARA5uHZODs/d
ke2FY3Tej4xJYDdfb9qaIkFwrCV40VPpGuJvOyZ1rxvNNmrK/7jTpVCDTdKHuZfAg4MyepgYe6ys
7q8gEn18wUWNhX0bZGo6NB5wQKhH8YqoQPQZwD5Jsb95zGdJ/pVRVExvPpahdi50WzA+/VFqNHKe
JhfoU0hiehPbJWnGSi8iyqeV6b/2cS45RtT52bR/BiyVZ2XdfSILqtgo5SSYtzpB9iPoaoEg2tyA
OKg+IWTWp4V/jUVytfsWDtJovqMRc70DGqL53d+xonF1+8Zw3zZAyindJ1DmqKRo/p8qC4/ah2sI
6q64iy58CjuUyiNK7IfDfI2OogC8fjhhBqbYu3Hdpfh5U5wySiR7IeSIV+asWAeEr0gFeO2gh76Q
CdIxQYm8GGAC5nlZFeeB1WaeoQErkUoLqh95teKLHViHewWl++kisW27UP/kUoLXacwkagbg0QT6
QX6wrX8XZ2eR961/5zPqGPKM20/mCxbi8vtzC1Mrw6SoD+pS4jTkW+uZwLbUutZRsaY+OMvq7upM
7fmqnITiTOKKeW9guBEShzCeT4S1OTtYxEjXGD24Sv/aCrDZBWJlWbP7m9QxqjX5MhNoXNj3Mwrw
RtKKC6zVc+6TLU+HP28Cmzlsto6BtoiLeripEbWDOGwvsBjfshuHLW+/fBiOOWTQk4PKBC9g18Cc
FPx4hTOJGHgv3evm3kwNzPwpZQDESS4594mynZLGQCSyt0Ctt7O6WwXLwpBx8AB16oNpUhqGd/3T
Kt6lkuKLLb1TwssnvXKoenjDisLeVU0aFpNa1W43scxhIKi1JYz4iG/f6eIzYn0kcJuuY/dFImAn
miK/OuMpO7XRyKX1uqsqcPBt6Xkr21is2LhwT/juVSwA+h9AbfTU5QJmj4vR+pjfc1p+oacBELBJ
yq6VaKEMZXihUvoipIXtIZFRXkSzYdFNWDulG9r/2QXf6l93frq5DLUWSyHKLIEE8lDzyae1olvg
CaT+hkOSYVPifdS6VQeh4C70+xTT5QefUy36pB5qIlFMY05LceosuU6aCgKfqnB+77j3Nl06Bp7D
vVOHdBXPrINz0dYIYFQMuH18+Wnvd8kqkktQdP1jctwUv71PYSG2ALp2dzHrVBO10ZFz5whU0Ktm
x+zC7Rsc8kmQvr4JUE3FStx5mDUYE7jNp4j5dlXvZR+cBHDokxkFrb75Pod20z0Q0wu+SGlCGR4y
F33UhmIE2PDN24dn9rhET5RW/MPrKry4D9oiMoh8oBWmCO1dSCajv9Emv84wkZRtgZpHBtBT5/bq
qeAINqsz/fgyKyT+9i5u0MzYs5yxDzgxbzQU3lOcOHlCFlV4dMBBLXQTF4GYXoqk+TKRrJgCBXxC
ETkEshLsvXkbvAqjV5F24QQzMoSz7/WcQgK3x1TeuDe2nfZZI3wug8WGSc4B6hWvkNuPxCkjijLY
4udTsxoIJKoxWq/g+AAQbX+XvVYDgBVREHHghVEiD22MyEFSJsialkcysiNQ+SzzdZv1KvO5CgFo
YDeqG9Eo/6Iw6sBc1PSQW8W27fhfSVezCxN1rKOI7kr6Kp9pI/edzSaaened0OQPXQA9rnFv7AmY
aw7CzFde1/gLu8+H5WUi2lYQJQ7e0FC4Eb/7uXMtRdHMY3/QC5L2uXVtRxrg39FQUFqTDcDL9jrM
ruBnkPSdoq/MUU0T03z2vzKCM+z9GLA3SAakvDU20L1ufs8928Bw+f+wiZv88lkDG5KyA65PePgZ
J2KJJl4rghKfxyDorHSxDJ0sdowSwHEw5cIxtQ8KknPPVIA2vdUv7UDFsdBm8taWGuUGTnMVtp9T
UWBfYo+twoISw6VGAeeS3LPub45Wk51FGyh118Q/Ac00z3FOj8ibwuzCqv+H9nODaCQHz9O7MaMg
SZvzFJlCR8r0nufw88VoKXnsu+gHH3ts/Z6VoHERGgZ2Cv/HVjLG1TJsEc3wjUC0Dju3grzymP1d
LtE1D8A+mqg+eKzDqxeVMrsqK75Kg6kUJJYu6Bk7+8V8/sea0LNUS+j+SWUQfWm1zVkehkakMr65
VxaQYSYXUlltlIm3998ER16inQK7a1s7zz0e9DYY4a+HjRzEsf2ZzLDVXA5frQL9zjDiIiVqoaO2
/bbtGAu8XkS2STAcPYp8d2VDAANT54OmGm6+cYWq0rLukP3rWYoCDxfTG+MDTHvk962llVnAsKyg
wj1yNkbkieHssGqQbfuZd3B61YKNqL+k6lPVbiRIclyx3G+BVnI79Lz6xW9MeADAdaizJBm547oa
0ASXeY0ebDji+QfRmquxDFxqAkMXxJ2VV3eO7XjgfIWU67lPwS615k1BLARHDhUomuwGa9Y+zU95
iEy53sJHMyuSJX/2BAQhs0yOuyS71NXpuChMzsrXXDc0QhyFs0MNauySu3CsKQ+Yci4MhMAhKc+K
8ZPucP2HhpRBSB8lI5zdGz+Y7ZOu7Ht63tRraLeNhVKuJF2Ps1uOzD98McReKJ1aWtCAKnOcCMqH
QfxqNnjSHrnHq/FSIPbxATc6reD0pa4rWTmbqoa0UVahCQIVG+XuYeW1v2G0OJmuIMskIb/eNLJt
UC98oOmTScXzQRoRJjcDGtWUH2iQGgJdM6BQwfq65RS609H+1FGDuNQnDQaL+qr/2qOiN+QTJQvF
3xuPsIBh82SxGtgr6cNoK5qhRrg42u5xaBfqJeuBYBYXXpeY13SclSUFFgaX4P0Gy1ENGhwiSZkx
SkRn3TfnjCNQqi4d9Bm8t5m1ZBXZM4WgPRir8JVFtjaTAb/UDMyq8Le7uRbr4O76gUkGXlzkzbqg
VBdzYRuRN6IvQSYeXK6GXCvPbi5Cppx4hFs6G6AAU67UiUTWnEgdFi0FvgmDvU+brljlQxbIXopc
xcW0JXkCNFTJl12hD31w9UtIkzzL9raaEw/8pQPtPunrczEntH7w/1bGULbXjsOVsC5BUP8TdxuT
JuSl/wsIP/PtV/aMqsaEc1JBkIlFkD+tXeLnbK8hm9myZC4RC1XU/sqfAlOQEzK8r90dFM32IeBN
/Vh2Xtn8ZLlibuGrtdCzqBLo8s1oQhPzDOVY+l8XkoU93j/+zHxRYxZTHKXs1oABPDoClrxvAJCi
/DVTzvZOXeUD39TewrhBI0k6cv7yHERSnohUeBpSlXObCWX/Xekg7rxmO3/5Srfb6kX6M4FyDs4W
1sXUAgysiVX+dGgH2PxK7Vpj25dP/2SfAaSoHn51LlESqfLYa7DO7XVssu+oHMxqbmQdj63jaEVb
zC6JD0rr0aBgCBAm1B2tVraMml2JKJDiPFZiGrXRXok7fu+hmxapj3iFHPaIqJjFkuDro8+QG/MQ
ohX3xz75wKcF/xxZAMgT8MQ0ZUeYz37vlwunCkCjHsuJJq7U1nKfJFPSgiJ1RZOQV7I1QJhAIUIz
taG11WwQcmviyZpbIQHxBGinQ6yb5j/JinX7eqLJLLkfmydDH3IR5zU6rJZH+M/xktyhZzVfTGnY
ikIOtmCpMUBLwaXFFpef6IBobHVI4OJmb1XQwGlhAgkIPJcn7G2/7NTLHp0O6Sgjghb6elMq+Yjr
muFMvsJnvJV/9EqLqEm9qvz8lI7Mt0al6vb10qOvnySJnJSs6aAs4/40dJYXZSWFf+yjtBE/Cd0W
yrFmWZ13G3KAgL7E2dfTnLo6PKJoIRFf3fB+IyutUT7wngHVUv7reTXYH0A1Kzff8edoMVE7LWlK
tN4oYU0Cua5n6+USeV3vvO+ahk5TnCxQIWx07OozkMYvSj9tE3+E63b7yxsfsIcBTJ9zozUoTtlI
TvqqDVcY0OT7PpQMcRjcRLXB8HF4rT5UwWiA+hZsuhLyCKc86HJ/dOKZOTR2uWGrFe3PwnkY8aZ9
zxy/4VsiOg0h/bm8Ynrja+f32quOVWzxtNNs51SMWlR/orlf8OYq49c5sAG2ue4Ap6wmCc/6kssD
b+tBP34Q87M/d30f11FBwFScZWu6w/yBzNbHJ4MnAE+dmSm2yh1yZqHvm68rY2VC8gxlTke34xJO
E637g93oSxNtUdaggiXE+YSwoSEcgafIIWClAcoQu4KeTKqLoLtaN4wQXtvOhfc2MiD0v4P1sjDH
PkQzcnd/OUcBIDLzIWWYTsFLQShvDY63QTINcAdRq/94v5mQoUkERsbg6c64OswmSKpl90Yw1PH+
fXRg7Kxw59YiKCyVkG1lzAaHnU9T85TtqgKXnsuJtXVgzpDL76moPYWSchoOXF3EblY9xLwr3pYG
NLo/wZsi4uxe9TDqE4zff6YQm9XozPqu6Pt2uTTQQ4S+i4iE/fxZnht1/+cl0GNoc1P/B6xI8lHR
cQlVFFMICvqESmpJa2X3eThXSHHsXvUzEeSQTYW5k2SFv3I5m4TIuD9KpuUcEIuS0DhMX1EiTfGU
w5HNwC6ACxuOnHAw/dK8zDTWCfeeV/rr3t8NjlDajrA1c+FRj4gjYu+fiva7yEWjxIArS9/YvJZQ
z4/0vZV+5VpEWSsuuLheYY/9rS2VBIEEXBdf13zwjlKCba/6Krv8anR77Vk1lFkPpelrPVRc6PJp
Ds+79bBVXFjxYRjwmcOe/NZsO6O49MZq0Jznr9u3dByAOvwl7j+8F4M4u0dVLVUY6ATnbssv6ZdR
u++QVOB5NR+E9VS4p1/ZApnlvjEPCrG7wT86voWQXOXpbgLwVlMwLpSa2l+BB0z3Oraiozdvfp5h
vgdkrp+J04wT3fon2I+30EwnnD1l0NHkIr2Czt0hqTv6QurWY+OjO7YWNvKWWuwuMQe/QJeDiwvj
8DyeBilU0pcnfrLbGL0DV8h2bIQ5b7uI7WqQNsZb0JJ2Yvhv5rekPgi+RfZzK1va+BEJnw6I0f7d
vfA2WzaOIUIwfYTIsPg5MvfIVMaRF/TjXy4/phg6x2jaIulGXFbmGXcapsJMZqrPfs+FGkBDjJlx
ENPYpkBNZ9ySFGLnWqpRJOZl/owfCTMm06Qf0jxGllS2KoJ+FrAzhSekAUAw08iNPTvvk9ml1nkP
3VQmT/qvF0V9hdoCBh9uOtJ1uPc12oTS9tfTqrM92X7kNegdupv3GQBP2PkYswdgSz4YX0OhQX+w
3N4P4wQ6jWkELmExuX6eX6p/5Fyw3F2n6wTnxNnjVTD83kzXEV01MaVf4PyeD+Ml07wZx97x0tzE
22x7mcIMUhyHwj8XyHzl13UyIE680OikuaBZ7vdby1oW1p0Uic7twKhZ5TApnuD3+liavA0Pt1HA
TkTwE8a1TTotJNOGEb7aE7jWG9eRThqFemLkcUoHpM2KIRX5WHjWjnNFvxxU8P6bbjCsDLtNdeZB
Lzdtdfql+peUwEirIsNUkrcMKRNk2pdmwHV2wpw5JU5YladFdahm/my4jzJGqIrTReK5s+pDpOgA
mMqXGy3ZgyPzovWpLZPliLpAeEeG2q+m9QoOLCJX6EK4p5/sZQRgQzWR8kxT3pxwX2fXofJpaF9F
etG/b8NZoKQwVcw23ebQ0i8tcqclCFgSBwbcxC1BC3F7k+GH28w1kIT3puXjP7C87J+/d/tMt7XP
SQCqhMCj+UF5ctiShQUzKawxQKxVSBzE+kC2N16LfOm53OQM8PGJwasMAwj1ZlEVgRLDKbSe59zM
w3+vbmJZ5hxzPSNjCVHrXntpLt0CxUXCQdZRZOIZLi34BpFzYlYxa0/vrQIkKXUD2jEcdxgjUYz7
UxxeAkh0aPYoOOJDRlpGy9j7l5a23dE87HLsmPmUp3cGRPanfZ6c/KMD/+izVlWK3xT+r37i+l1c
H9T4kqJC+zCxerRDPmb1euNXAX1jMaQ0G0jDLb/ShlI+va5yXr/K7rx9ruq6Y0kzSZx8/dxmiEAv
wiHMYcpm5sgChh1cHU7rGSyV8AL+g7d525eoQqidmt1ds22V27s6botkrrnC6on3qh1CvRajMXsX
3o/+HaapqlJjqyeBQc8ElDEDVORagqJQ7pxa20JTF5gnwPM/jmyXz93/0mJ9DU28noc70yeEL34b
+eVtpCr/jNVHqn0qcZsr7kM8pji965VYzOj2Sxpo0POfPBDWJv99P0BOIXwsuXnzDUuOQPN43nh2
tqtjH2OgiRwN6vySxJ4qYqW9lpxk3CBDonOvnsOjFXh4qUKp7T7DqrhBH456dw8RRrB0tTd1sfwC
mUuo29PmeqibaSX39CzpRMkH4MpxJcP6j4S8NSfbf6VJ0n+tgC1bCjwFYk1mfXnFK/IXakF0+wMz
7gOX18HOyJm5rQxzKKNts5sX/QugrYP4j9ruqIAxf27FWZSte/LcQcr9I1i5GQWOrzkWSniGNpWv
yWwM8QfjcDBZU+Xujl9RQOiKS5BdYIw/AmC9WCZ2u6etVsFaC3StcEMINymdMyX1qmkImPQ75gxl
5Kl7KgaKoc+IUR8iFijjBSpS14Ihz6of1ZY1Tb/sBkJcqs10cU0qULpMbAADxwrEOZZi8h9e/E9R
2puj/p0VCS/Wbs3KVPZ8lJqn+ScTLpTZ2pTMzwGUuD/j5pXkHItDob6je9lYrMYeUxcJnuYsVXCr
SUpmL6scG9Sv3EayIO/uZIACHs396SAxL2DugInyFLZnqHzXd+7OowAYfErtpnizmKLM51ZpRYd/
i6VMTDckZl3PAcc9hoQLL4FVz23uYeTbKN+1SKYzS47Fj3owCH7PWtDlwPy/d3tSwHfd7rPvgOwG
9+Q1ElDINdDWPCiK7NbFNoDeuWrDzMyR/zAnzo6P0STPpgEUiuqFCGNo4q7PrAappr0GAX2XGlKj
WXte5/RnJ1gC4wyRjeR+sFNfFzD47lXjvS7QOJl9H04Rnfly83Bz5unbcblf1ZjGfSa0ZrLr4QSR
V8Ptd6rvdklMLvx2RKAO1dU4nRBcK5MuaK19BCPL2Y2h39IS2S1gfDxFOQfDyPZRltPA/MhjszRZ
yjhhfZTeAeXZM064Ui4Y2gZg/ta1GSiu5O7Bu8cCwipC83tOAfpA8lfoiJ3nB+9O1QyEPO0hqFCu
wDutHgqL3Xya6FfjwoV++tI53d8ix3eBi1s2AXpRipQAYJsoDLSBDhQeyriJUACQx1RpIs86BBHH
5Ce0rfFU9b+BH4EMDxWhKyaZMwlUE5GsUp3Ycbr/rRpGz2jBNAUob2keQmdtpY6enHxC5PmQ5tKE
jskBlGrhAcYS+ZF17S/KBQ5H6FPut0ivj2fau1v7b04RWltCM1F/NPSKqGamqSPzqAZOsa6f3qaX
NlntN8sqHDFXUEJ44q9oVPMqOsfo/g0Zi7cZgXSG9T1eP8kQ0aG5GdYpEGSctexwFcxl7JF366K8
xbZX9tRtWWEr+MUiogq0ujlwoT9qN20lTp5UAjJDG8vJKaHfL9inbUhyxbgVWn3JSouKjZBG+Z6h
MXHZ/bVPlu1IusmJ+a8hT7QUSV3VbvikTQ4fzvxJ1IQG8d2E2D8I6lRrJw8omRzuVCwEqkZb5VTj
v4l+3tpArYouQR2obqOvJyJIq44gTSqqQ424ofQhajaZ0/KamYJdj1Tvypod/vPIdIsppq+e81Ov
lMfL7+uofOYnVKWaa8dWMxcj0zoLLKWxiCLZnaVasyd3C3kivIplKOQPQwTZcuLL7wVpKn7zJ67U
7nOJIfrUyksAqXqQ6Uai69TrjSG6QX4a8EdIIGAb8ZQuWTg+McJTtcrS5uml4ET7K75Wj27Tx2Pg
GO0HA06ZEMgJFMTLr6F9ezV+puBeisod4JG+97VVvqP0JrPVirQClnt58l2uXiYMzIWQN3XNjD8H
HnKTfw/VeXZI5TEZVvWmMsM4GojLu92ypHDrb82k7r2n+8c0s02Sn5gRkZEuT7D/p+3u5opVwu14
2rp0st0lJa0N4VUv5x7fFVpx1tbXg60g+0K1BAdCrvdDT4KlCPXV26Pt4J+lSkhHuSRNFkwAQuWX
F+8m5mWpmpbcZUxyl2Bmtdza5gfV8g4BVWyf7ZN5pcdBsviK0ecvfTDrgsl6wia+DkJSoBJo6HMb
UOHzNPRaoknUsZ7Q6DCD+jXrHrqt33a8lVpBV9ASSyHp4neEjj3KY523ZBUXpqDk0qpXoxtAHfEA
5Ft4vujFZ6oPE9R++xvMj6Q8gZEJkRZ6yYBneddFcb7ot34bP7IO2ocS0n/xW/oi9Q1M//2P7Jo1
7ohgseqF/jxJ3ojyrEO5iTn57+jQeGArYDJTGe15JvI/KPEDPDfPE9uhyYRWoPoLeoHRLcOn2jeh
9BVuwbVSo4tDwNJjWmkIRonnH62MdIzbALrj8EHa+fFl4PYXJQY/0PIJapbIlrT66PcNly2VLpwc
Ynq1E2hIVjF4UsmPCdaY3e13jT9km6p2VAJWjgB+5ag4XqWIzSNOQ9eQlo3R/ILWAlgWBI642YPD
C+Urpte9/PhZFdzl6WsRciISh811LDveD9Obx3ExCJKB4/91QwAVs1apHO31dEMcqoGnNfxgZGCR
vxeRJSvS7uttVtf8hmUQNYgBO02KzYVKKZ82INuXVQP4DJAjkjTHBJbYgEgW4RuQX5tqi8XlcIJ0
5WydK/1OTt3WzLEwZKzjEx+LUIe4LdJNCuTIgvMn2NdTesADPURGb2KXNd0UdA0snxrHZubzmRZT
doGGASEBSPzYHrxMNAnJPzZCAXCylcmVp2u42S4m08PIGljV01B/FZnP/CfM2mHgYWEkGYolWf7c
LM/MHdPRkiX//1+EF6XBM60PkM3LW1hy5BRZkf4znT8OtajdFpbx/qXjiV928nWyUQe+Y9ZzJiky
RAdKD9hfRIDhRmD7K7XPhigU6DU19t2QCPbeVR77/Jw/KpUOe3KChWfSUAVx0L8RoDxUaDO/Sho1
fbW0TocyB4jGh4SJhNbps1ZjZtweP7vykc6eYwRJtkYHY1bx5z1QsqGJwVngmp09ZePZKuiR2tth
HLuR0xfIczoqjnzlkmR8haoFoUyuOdnCNNOK1dLOFhJx3sEUWwKOAGupWanAZQleHbgH0yx9+SLB
ISn6Ws2IO2F8gQio703pmu+tGhCf0mCGrSfVbloZ2iFViyQyk612i/Fa6w5KmwzWYMObBb2wG2JC
0noqB4dzlubwt3ivs7EN3Tqm9eJcYUAktKmpb1XCo/mG+U76CCAs61GSdAOnK+21ZoPClfTuPA3Z
zDqgqg80qp9MvEK5I8Qnkip++ByT9dPgPGQ2FLbJ+9QuVYjE8p6I46tFFnPrxlRJhlncbUGjYw+C
/YTAqWjgr9t00s3P5Uin6W4pUULxPzwP95ToU8chsJ9oz059J4z0P6KPd4aJSMzlv7aCLWKrp1lb
DBAKZPNA89oaOM5s1eAhatHet6DFxSFAGoqoBinEoQlzvenl3JGppo7x2rLseOaBWJjB2iF6Z+Rz
+wu/GZTXM2ylorW7QvnBvxi06YLcuZB7bH7v5BuEVN6QtmpoiyoZ2NJyjvPsBfLAoBaqewvontKr
Ji2iFO+wfTK2+if3/BlAEhl/J9ynrKh61RkL68SZHsfXAaxv7Edmra8NgzTLcW01duaJjwYzCbEO
Gv/fkX9ptlUMiXoEdXilHg3N8i248xk0QepCwOoxbNFGrV8GctYdqVqO+iBwBCALUzJYiRkyEBYn
SNvA1YPI2uSIpIAdiUCXPqUU+h+t/MCLY1BFUupi8QorRgJJf43jqkv3EAJkPklf23zI9T+LharD
2Snz7TYiyRCoQsS2fA3vtcsV3HpnGoceF2v/LkinkSfZRyHhh1XLZu0+vOP3tMW5JQJgTAnnHjDh
odjmZRjXcrleOyF6omLF8x86Heaq0CaYyLQDsLN2A0QIcE6lBKwdW6ebqk80sTf2od5JmZ4UyXGo
RHTG78CL6VHfpXGO1M0r3s6GDPIoUSRwghrAS2zQze8gmaxTijEW77I10yu0sEbNN/WcWwx71X5x
9slq0DO2EwkOgAH0mqqKozQxQoAqoF7Zza4/Orb4IVozZx2GJhxnnsjL5sQordfp57hOZyaFDk4m
D33w8y6NnDYMvrnhX5W4Eg/5y7iNA5JyvBMF1pn0cAPqVjmczHRmRogK9m6ujlVq434hyF/hKJSg
bfQIycYVVmtUPCmsCc/Ipd/UgZX93bHCWh3syHG6TN7SwAWmN+Yt8rZxJJaMiqnfz+jEviFWofNq
5qtRSWfNmU/bReVmGFgiNeEYHCq6Qv5GQHtncp81H4L90fFPvkxxNlTqSLOkjZVKawCPYkUSiY6Y
NhXSp/O2eZaSj3Fe5oqS/Tv7dAY9iETkr46uhoWv0wbHofA/0SAf0Y8ey0MT1D/gNh5awWbw11lG
sjNRdnsNEi5odH7brqbu7rYMhINWcNYBjpkXM50HCPbW/6AiUCRH9EyGR5V8AQIQHFmW1vi9naEO
GtuNBAeyQXzeHpu1ObnWCf5B91z9y5Y2FV0DNR+0wZ4gZzNOHo1UnUx7f1DGDDv+33IPhIec6wU6
ggg7/hdhG1hTqdC71HdSzh1JM4cAiVv8FS/D4WGkeAj2r07yLytmLiBbhRWbE8D8W4IsMSelwNhw
vyotr/IQNGg9+Kv6yQkkXAvh91ByIdD1tV0XKL3ahRge5b4DsWp+CvcccoAdQc9Yqn+ttfop5E2g
4FVSdwj/KTucK2ndzRiFAp8u/K/e7du1utxrod0i0SaZcxpiPImS7cLCXCFrj+Mzqspdkwm3xYIz
Yc6nXF7VZS1gRvfi4s+xOT7n66gybIWY6QVVnyUP9P7w40gSxhcWcddFSTSdxTCabXExxUKVszD8
9bzbswKdrS5/gMAuKXL2a7RPCxh8yIz+Vp8Of8yU88n+fEkfJAhRH/a0y+Pr8fD6YgBH/vjalxph
r4btSStwkYwGXHefOOkbHmbCFTNH7tOk1Y5bW3VJFBrxYXLzUSC/FQ002sgdr8DWMgeuyG3Ptehr
rAnq2hWQaVcWQ/I4dAgVPF4n2+/EoQxruM10Ge8okupMbJpBafcbRSI7Fxi2hbpcqOPKFdnQNfWU
mq5WAaWI+9MpRIAH7IdZoFc3GE/2rtZMnhJLyr9UBpNBwlbjEuSL2npWxfgiQvgNPV8egBHIGs4r
DgO9VYi2QMJAkWrPxJtre6piIgdHkmuwfeyJ/BDEgNNds9mCjgQaeK/1FK5NyR85kz1UWlvfANcZ
rcc7una6oOvfFJRdEqY5EEFT9llIDyLt2vTZJi51j5bAHaeyeuLsX3CH3t3mitT2S5wykm2JN7eA
DRXQwDR+hf0fcnThQEKJXE/VGmCVgKIBNMeEEcSPYlTmGNxoqMxC7A0KKmVOZQmzFew2wLMi5iUM
0apVcbRU8Xbr95AXvlaQrr91bEG5mJJHMyMJCjly3O+bC+5uCYXLirBPeOzsreOb+tAEX7xXFUjT
Nr0j3HeW1z06vWrfGTNw6mSjDHklRHwqbzHkg+JdzXRrXRteRl0RoWGTAs7QlkmknJRip3KkDb9e
iTbmsQM2asE7I5fKO8OZFWS5US5e85hd3nKt2lLbuZdHVY7IxB5bt0jzMlrRPM410mSz0YIOpGUt
yfxTFr0qscCH9U5AgfqbsXaZtS/nCibYilkVVqT38G/3k3guZJexIZJzO05t77/b6e/qFtYX+gGa
dkdnS0y7HFtm1HVq13+IZ75mOI5o0mN4+MT0a0EXjK9QivTawuUH5FiqUBrUMqjF9pfRa9Zv7Q6i
xX9EiD2JffiJOz3p02SQm0mDn8rD4G2g2F7eUnn9vpmr/pLhjt/nNyohdTODoVHPAAMrZvRnj4S1
43V6z62hEBjrAnB7nFpoflm8MDWk5Tv5FuOlW7/y/ywPpv5ZDsejw9SLHXV0GYb6IKvOSC7UoWLt
j6uiVJQVIfQWTNPtImXJW/oxZ9PEJqcQCz6FQr6NIQxrAC1KNpBWYOJmDHGxh6J2K41ESea21XMW
Ere7eH6HWLhq5y4osYLCXMe9yatHhe1F3JUN/j/8OE077ofkfnxVYm40CUWffoEhoFmJLQkNVoPd
XfEKR7XulTexouH5sNbuNgXHWHQf0ENwCYApmWEq5XpNKIW8wYwf/LyEEbn+Nm33FxUr1QrZpBSG
facB5diMeLUu2FEfv+usg37ue2Vpap48hcgnRfWnjz0/tlDqD5M5Aq+ycAEoHnbzGS7yTaz9Ff/3
8bDBcD0pVRHCWI5GG+LmDgWz0U9UM9bOvd2z0xy4PX6J2fVobewuVbcONX1Da9UOLZ/uPmFwlm4c
WzQ6JjdI8QThu0c8KAZO6KrqlHFSnG/gXM4NdgwLyZSz3LcGML9qFMqyxFuu6fPEpm4fcIrz/G5o
mY3PfcQIAgWoGSP/gPtKVPJaMn9xSPnlb2vvAW5KiByDdKjKNFZ6gGSJkWSzxrOb/7dkK2kSbQRa
Ma+Y4awm+KwxTBOzEX41m1LuE2YL43jU9/xg910RIu07Rk6tih+p9z8shmOEyIhMKfz9iabObRy9
d5OktbfGdih77PW228RKqX/rykHAvc3RAFSNLYBxPQkZltvYXkBVoEg8hrnFmYAWujySBP1DKAFr
k/J4swILaO8zJ4niIsIfYt6BB3arLHsmv39SAyTkqtnCwGNUvurMhtCmK5PIZP7HjDrMLnjyuy5B
9I0yV5BzgVzRTOyD6os3/CJjzaW+Qj4LmzOaQZR+dXD4Mg2Gs9lI9LOcgOgbv9WzGzrrVvP5hVLG
YSSOTRjBv8T/SmdAHgr9LgdQs4U4k5jPhzuxSc7sYramez+cgVRx1lYM2My7qhuVYTyDx5vZ3Geg
C5NRL6wGgPL8jEwHth05bzUhVrhA230/cqoa4WlFSZ8zIBF+0QtvFESgczXv8JnaExVoOiwvLyp/
1cAgmVN3zjenrrBNK9b4NUndwZbxGiKYOvzpVdO0yKbAlwwHGHCdKKxCjM86yMDlT1t5WzYUJN0o
c1kGEhgVSFM9LTxJIaKaaKrPJWTQe0f/qq46qsVBkknlESKtHFbry7CSXB074fAGzJTvhAp+2QgQ
ZH0ZLual7RJfU2FGDAQzCEY/bRQ+PFiDQ0CIg6PLwjp85N6GBj6PfYhnsp8NX68wgpUClCys4esZ
hrN1YocLjm2hdjDj74lwLqsdxHf/0TMHXKInAcfD8Mc4x6a1bLZInL18jg+Cr/JMclzCJ/eLfubb
/hofOEf1LHKzZ8W7j86GLpN47mfNE4GNH5QYslL1det1kn1PcFYKR32uOgnIca5p6WL3x6g+nc6S
mI0gNL2w5cs7XOtjxZ5bv1RWikjUMXBhJ3rcRrHtVKa85FuqIr0za8lJNNv8X0ZctGu2jCRdowxh
zeWu1ucNPQz+RAHSM4l63FQaqh02CyH83uyNLsLe3VhyDJ4XtkdkpPxirng3yYvrT03QsVkANHb1
Gzs2blNnMgQ1YjbQOLEBvB8YS8KTuvYhhIRKHF8v9IpENbgfImNWbvB5PeXeyd97damrrNnEVgTR
41LadsEiOBak/bhd/Zt/k3ZF+XpraVT3B5ViZprh8WwEOK5EQcF18ZsBa047d7B6geQvfqpiNNXq
DzP7bPaogjup07FwuA7w3DmToctBkbG6xn71mUGeXtOvvp5/E9JEgWgZCMgt4SjO/tpMXvz6pHX4
kr+B+RPBXV9DBHyK64nOenhpVxUCio59OPIkQUaVnTWh8gIjdM5n8dtLIKv8bWuiGyZb/6aOzmom
yMow9hTs6Ydtx0IzfgOeNsPmFBlsCv90WOtECBin0mhcAwUyrT6SihreOrS3pyJjOAvjec6OgBJW
2G9w2KJY4HpNWvANV2FpPq3d7bfh2kmzhm3xTkAZcVxK0fmWSWdoCg/OyRMlE/t0ZO3qEt4qJjWe
fYBDi1x8MjbWCBr5y+ZOkhxrXh/nJFARJcRkZ+bBsK4CjJ1puj1zW/4eNMW7AjO6mVH06AoSvpd7
QhgZyRCnygk1DCm6mCN/fcGpljtVMXxDWw6TaYh8Ahgg7QZC9JKdSsvHZj/vg5KKhHr+PYBytnFp
By91HhuVR9L+rBh/Fm9z0ebnZkVbyAEKucgyCurCYdaXgZdifzjXEEYIF4P2mkADa/xjTqCfGMVt
AlJLm5CntLXvWqWdel2hxoWP5EhNo78PRTFWtxcH21RdOdpK/pr9JOyLwj0jvA+KPSUTWLiY1CEn
s+hqBPPXR2a91tzs9SosiEpUVhprz82tsw5s3Q8YtACPfsf9spLYhC/yGe7W8sWuNf7PEy79Puud
l9lFLHa2TxJROtAGgE+kMCOYMwCBkrY5BuB5w9WwYtGGRHjsJKbq3aIdJyDJxHnVWNE3vlVNTUBz
Pq1daZbLek4PP+4Npe99/X2DpfYI+sH3FY6KyCJ7HsHLyw4MAHWgPXupLzChr4aa4OSTZ/kGAx8t
SQVVAGw0xuhWc4lqEtWrSVIfY92IQslgMj2Soho8ZURpf7R4dLE4P8UEgZuTWpF4ol2ZAogfcgXQ
y/lQ2ohPDLo58pB4YHD+zp1TGVP30Fhw5B4iAlxL3lGo2oHpo/jgpnG04Cl1CrULEs2OzYHO01Vj
1+DjsMJLZA96LSTR2tLkKMI40QAuL/C+/SowqGppnLCS6l+vAR9TTs+Fhx+VrBGB0Lm1sJKyLcbU
BvRFe9SIDotKy2Z94KkN3qwuCv5DyeVYMSljWKRD65SeTTAFpMOrVfGRAAE+d3nsg+5r0ruWGPFP
zrjZ/QVK10b2egltt5DkY7P0O5c2XukWPX5zt6gHzreX0qBkG/gK01ViTn0V8UhqgLrZFahYdtPj
7TjRO6HkezePn4UHEyjb3NxObIh1oL/e1US+pOi7lIBbJ0rOVCAp/kzEHXlboj+4YscT17P9pKr2
lFLg6fLZm0OB076cz3SNgn7NfRYBb31jca8wO+XJs/uIRevL/rhOurUc1fnGFa3r+nr+NEx3SRhq
5RkwV6WcfiXid4PB/Y04zko4Fghqes0D38jDiKQoT6ZCQ05+pFd9zGdVVMnNV7vcaswqZs4I362f
MvZR1yEksHDuNWiuzS/XgONnei78ReaZ1qt4c/VgZs0XiWUlULaZJ+NrMsBlb/9FkchyUjZH/u6H
lFLN7wDN5jvDXcC1071duubYLM4Q/YPMBcjJ6/fllQuN+/6LA+vP0mNDREkP8Jc97s2SPsQ0O/iX
eEl5MwDv/XdQgqJ6Axqipk2S+YCknrNt6Pd4yZxHusRRasztaZY2ApBWOmOfn0WUcZrTGpC6/2/U
JtzkCglGNFSYNwfFLyUu8UUy5A3Nkf7OGBo6tXM3kCI5tYulx/6SxnrAyXFVAaWAhHXMUusOL4dh
+K48+HS6i5qSUWjpw7slpswfDXC4XSEVtBj4tTPHysHeBEwZpCcKtm5zjG7hWhl4T/9+dN6TmZVI
TSeiD5t32Pt4KmwQbQvxARqGLFjPI/hyVfTDjyLTP7G1PAkLVDKXOMAxYZt6b0E1lvamQ4rVU+oI
o3v3ilYOmyzaAM6kSgw8Z/EMvDin/BsrAer66W8qMak2hBDdUHggSe1Pz48y3zWMEulI2PKuIPzM
wfl3jCDoQQrwvTYZN8oWQASWmGNPGRJu1K8w8DKRq87cCawOzIGTVfX4j+DFVcSOTC5D+n/yOc3A
U2U3q790226bYlVTtzfos5DKpRFJLicAChjtxUGF13JzNc6MNvP3fjaLDCYGC02Ut91aal6EylbR
4T/P/j0K38KUaok7rASdZF2J35Tm4e5+jM0eJSeJsq+c9G+cDDhH9kwa2UKrWqX8XZ8TJevR5gQ9
U6/LNkhpIjHcugNdM5/VN6SL+lUPWHh7bzgwWibk7M4Mbi7909Wl1Q69JX/zgLTMhqPfyUIVvg3I
q0rkQ/3XtEkg6VPGqJXkyPUhKRjJoibTeq96H5Lq+zZHOpJhwXwAPPLi3EpiNDC18/vbQ2HNAn68
3rNCAjEhfb20iP5/AwjRwR2RRhQJjLmAIMddL1x66mCKi1rbyEuLdzjew6+EF+LNI0y092axKgu6
0HsHpdVE19oLFtqTiF0CKLhmuAwcPolqV6dKnQ3bBuwWDQIlkR3eK44m4fUJE6MuC8Y8PdsGrbmi
mrlm+xVhSgcltVWCeDu1JaTh2oxFuuPKJpTBG4EQSDqYBuqRdpUbuHWB2MQuZPJYTwOxYY4lLD80
Y3zZro6MPpHjEFdJt/YIaXNiUPRFkih0ivJ8zzBxawJtYiVANDf9HFe94cR6bEp4egclMBDVDN4C
PtukGmBXHXTg5sNxEbYboGyKTd8zfRJpQhTi5AtGLxEtpVcSVt/7pSjErDxoq7PK0N+kSjKeCZox
oJNDRAl8RZ/qlLXioUq1vEn5iktxe/KyapgZXKHxQxpjm2F/Tdk1FL573VX2ZE5Y2jc0cte3Gwtv
fsiPSSzdqtjriGNwyrBjSeAcPvSC4P0HG+q0vaqBHNa16IqF1qZx2Vy0Ku3ilnJNHBStnOHXUgIV
TIVPDZfG+l0NtFWFKhd3WOMTM+Xnc6nPdqqrZjhzJSE1tgKR80J/FgjfgMJpJZw9VcNKv9hDN1TH
40NZISBDNSeYcXNSPmCXO0CaWE7VUjZyhJr2x0b9s43EyE9DKVO1IKY92hPE3ee95o6pwJkKzJC/
yIqtNa5rdCkZcivkt0TnyQ539otLePHp9iQJfCMA0PUZcwSCcgbFwPlI22qeknVpBM8Z2aOOCC9Z
ycBdJtzQeoATcigeDoFK1IquvVHRw4hwEzxHGiP9PnK0rZuDjXdvBOjxTx7UdBnqHWZG7q3VRbxj
I8rixyTGc7RUo8+CpvJw296Z915tEps43N6+c3C8bI4gTOTaMCWW02SjoWnLtfs3dg0IupZr44B+
PVRIqSoBWZIN47OtFL3PVlQCGPb5Fya3xYHZBOIlFiDvcTafYZd+sW0Giwnx/71C5AVPV17MdiDb
X/QYkZUN7vkJkeIqexYtHyCCuNsI55KPwRfe0/0lyrPQhm/Aulm7ZFhGKRvFMPt+hgfDL6Djewxb
070NGWlNefxiq8BVFNfQyEbHX4/rGpa7hNJ3n1j6Op19dFznmJzvWuo4+VbZBuW/gN2v7B2gdynK
y8IynTEU3F0p/9vtUg0zxJGA6Iq388y5e3JjBmYNwWKQslOBTEy5+NbRzmpIkdsYPIRJyiZLuYL/
W+1h7Fsx4UQ+D44Ib4mWivaSulVH3ICsph7bm/opHFI4Qjp815Hf8SN50ofqUr5BHZ1BW3kBBV0Q
2JvHvZ56M7g4gxme8eTgCWuzJN6yyMomB1fN4WrgJ+qxSigOBtIWIX3wGDiBYJv94KvSRbuljVat
MxqNR22jyLjLyQ7qBJeme//lLbNa7J087zecjFW9mtPVCc5wBLPi1w7K3SCZzjCYh7YYRjBeTIfr
orP2zHv+rjE51ciKgvnEBBGnKVz8bKqC+uXCTlVngyEowCR6AJCxE8rxYRVFeT2LivrIQJCt6aEk
485KbdW3CRiHpv1xb/wmKQZtc1wEG4eJARJtB8SBnlW4T6F3aTZ1DtsDGvCK/8jzPqTVpOWlemIE
5UCfelZR+Oa0vxfh4E0wSwmdaX1d+HQOPQfySPqTWeiUtS5uMVvDRe23HCeQoP2NL6vq486Re6IC
ob2BtbQLmC5Yg9IqJs22YP/UzSpAl9cmdykzX/izJw0uKoOti5qquHmAsJvVjqJ+Euxc14+n2HOz
7/8dhl2G2VZZdp6LMJk0cMeE+PS1iXCFOfjmv6flPzzKEIhSz9PI2PVnyNkinHj+8R5eeqMrNDe5
zSeIbnvUOdhP9OFGtD94mbyGuRBDjPLaOJCI9wmdDisVRRdQ3SEf1qU5dIBxhLvXRCvHZwXyfaiS
WBUlz81y0uvkm89nTuvGO5d3xo22paYPIpmV2MIqxCIhBi7gWzbmrk+I25HXFHmrwCuv1SHqniwa
70bJQBDWpXtQ39dGLHmF35eSB6BWDMqhLox7xtEUHNedW8tCxCMDosmwEsJoN2sRmWQwrbCWQp+B
U63siW0sIl0UHM7bcjrgPGTa8AOeptz2THZqblnNIPeD1ENuakXlCU8g2noPnQa8I8QV7482FDOR
qwt/9eA1SEHfpwNcU338QlpuG7gC125/0e38uInI46MKvpsmkGg+NJrmfOFPEDq9GauFH1bX0Vbq
21tLsK43DwCKElESGANp52sX54Idh/zqyOtIhk/wkU2v+uI6i1joce+aQCiIYijzClFUug6h8cBh
xzlyprRd7YQL2gdTEcQsHGSxJIUYLWbxJYGXK7+tx5PQSYPPMXbQhAEaQO3jRWWK9Y/UFHuUbXzv
pL2IZZ/OzWyl7MgirInqRY+m5KFU6RW8Fwc8hNxHdO18tcBiE/6XIXle73PrvEkSdVQMgJPfOBKs
FGVYrKELbyvjbbAR0kPPGnCmwvuQ9E0zHrCtD7FRdu4/dnFySsoMjkok18sYmSFaAJqr09Kacg3+
qcQubYh6BeLx76k3Ews4Tzm7PTB+XTksOS49eJc3gt31nZEP0sZXCH3Kt+3qR/QS7hkek/pvS/vg
8WQXiD3FON7mVSHc5a5aqCV2i5WbvHXicpVlglh65RRVACPCSs2icxte7zKwkNkD+2aTAJWjV3vn
f0NFqZ7pvKrOUzTeOGFFRa1/b+H8Zh0hiYtCCnlUZMO+jmLb7jZEC6PrDr0Q5bD9UFcL3IVI7Tax
y71zRmmJmJ4x5293CJnSId3ac5RxUWX+j9SJ9aRViugQSMfXxb25a2aLeCE3ANAx5B08mL9K+SuL
EcppxPAkfPEOGwaOIe1RgGSVXP6w1wXRWE1Eevx3SgBnBSNppES3aCd4WNS8wmhrLVRYuKAXqXqe
2xZvg+kew01OZTorJ+gmXrwFT032AADYEBE0dqPXfymPrnNgkpUKMpngX6aWPvm00PANXTQMwZKK
loXUjIEb2Te/MAVs13zTbQwpppCUvqOZI14cRKfOOl4TQe06x0X51J2dGEo7AwkSxX9W9sNE/HTR
ChTI7IFWy4X2krlXbwUisQMok5GKyGPUnx4vZxUC8QfSrH+eQCcU4tVNqOAlt+6jRNdo+1xxQvIT
KZZaDvBSLXtpF8DCidBgNa7k+TxrrEdIoUvRKdbZZIsbazTBjknorTF34PKUNMwk8WaodH6fujeH
VcXMpLxuzoiSA1OdxlHGbULnhd5XkOuyJxQSZEdlnINKfMbtaJGTTJyo6HK54X61YieImIHwDW/e
BfsIe3uueMsDV3Cp6DLtX8u59J4SQER/pODYedqTzf49ZeebQ/nfVzn8eSV+w7rvXrr1U2sIgM5z
CELzSiGdTZjCFr1qmKZ2zP8MAVdUYKZU2dxeSBNgGLV0n6f+zUgOEd+UNxil/2LYr694kY2GDuuO
dW1RCj+QEesKaJy29Rtm0RKSzN6/b8Wz+NSEH4OzXV6pcgsq4Ka3aiNXH3rHG6S/DRqY4Fo4XOQ1
UVkgDXByCK/dEl+RorN2KLMED5ph/DKuYKPtexcyXOlpkbJdAE27vNCJrwxnl/KCwXKfwZwBH/sh
5OAPig9YH7mHhNHIr+RXCV8Uej3jovQB4Ky/FkgToE7h5+NsamxXA/YI35FxIrttdKuHYRM111Li
bQsgl0NmOj5DBET6yHXe85YhfpVDvfyczKMMLgbNTO7PUJizwA5IeZHCruK8aM3NFtKiSi/TN0jN
wKWV/ZmZ/uyusTMCDuMMUhP5gKCITLarP5x5j/29Euf+yve7n+CZzYd3ArhAE4S0gP7ksf9mNyDf
4VxKtJA/nVKkr/dly3+qu27mRm/HTarPQTe59zi6Ld8RhB4M3snkPjK3qGpbu+MHalQPOPEDRudZ
1tXEtYru1yFMHds1d2Q7X2oMmJ7IELb6X8U+IMEr1cvEgyHUZleWSXUomM+5abFSZJKmfYqLDCVZ
KfLrec3vqc9Cb54I5vkfSsZMcMZHD3B1ubitslndzwzs9wa5QnddC4ZQ8cGEL+KnpndDspv9CeIT
e6NNqCmVcnVzG5HjhHQfcNQ8d0O3/UEp0qnci9mS8+Uo1Li6s4066UeoB0XqPFxm1v/clhecc361
H/tqaCcPQ5J+t+j81IYX2exDAQRYK+8CeIN+gQD198UK+lrsCB+Dyz+qrtIUtP0Y2B4ptJmxjkYn
p2XvYf+ejiqQzUBpDT9RBOemzN39hs1x8pVQcxCKFd4wsO+TDyROwoz8bQNF/wkpqTwyqWRImKxr
XW/F/5LtsxME1r1WP37ey7Zj6VAeVm0QaZxyPwR4KEuMfztCXxgTlRLkFNO6LhIK9MrCOI9tGQaX
ldAJRUOMFnPLuh6Gx4eppJZWkmT9NAWDhoyFxa8GwE0EJhjJ3azcn4KdqVu6DyD0dHGTN0ID5jP+
lpEXaC4cspBF3lSXk186yL9hLl3Ss8gQnCAFER6Pq3QfrqxdRcKbSJFamfmLm2t7NsipP5eHHPzg
xL9LtlAkOuSMB2776z1gRwXkpTmiEWBqd8ppBLaDiF9CYT+VU9PCC+8g3hclw4oINmZP7vFp6ir9
Yr9SwyaalGQZkyYfe3d75vJyYDbBdlTad/mp9O6Wl/lqir7deCV8G/cniAUJ56FLxiAtmdY4AFx+
xAt6ihQTfuKt18V8dx87TS/YOXfv8QRRhjydvz5mzCApvDkBk85RpfUep64lgmUwndEf/Y8XUbCz
V+sqzim0MfZYIrDkaXdyV8XLir7I4QcYvctSuskPHZ84HBOrl52BPYWaBwxkqF0B8M4TDeMIWMhe
uleygJXlPnzlLFy4wDc/xDKh4Esm3Lz8lgXv1p+ZFwYpxG+dCjJBERkfUvLQbxupRNdT9h53JDTJ
lU7tF5f3We1hHqxsSYDfN64OrdQSj1g5eqkccD/90kZB2zKEmOnQwOyq1HgbCzBL87S6/RyLw/7x
VtzmiLzpJ5kt3nbZNctR3S0EHLs3lzPe8a30IvjKIk1JlOZgwvs8Az4iYzGUYWBnVqqD0DRYfMsR
QTE3McTnJtyZWR7x4hO7W0FmDpkYKqg9eajuVEmwovmM++Pi6ywhAVa1V7rGeGjanBI7raZeZtqX
qE7peXh185yDZxyeyhFfZZn91kI0Sylu7UfBGg+tEf7uQ8sfti3F6ZmA4Md8YW8HOQIK+mRvaK3Q
+BDnA53G54GV4OBxdJXPDOuaBGW6Ew+kBfC8hLb/+EWxRIfsHr+TbVUg8v4CGgd2YpcuVckfDtdY
RiH2IBJm33G9UTrJkM/zGVtlTsT0an9OzOhdNji18chYu7YBIxsdHxaMbwaeJ3BQcUhkhUi0kD86
Jx6ZFvlaPnvsSy3AYHJxb3z2RApXA9Y3/vfTYXH3Qo5l/pSzRuEPGaPc4S+sM1gY4Y7wQCrXdCx0
0VFGVIc/5RMW+M4E6C/UFri07y2QxHvyVpvQDXBZegBPdrPxdf+vuzKWmiu+Q0WVk4uo9rEsREGk
rGLsFIZZrUlv8CXJgE2HYBUhYYrfjpPE7uvkWFA51U+P26ThPg+w2wY3ytVWJnBZ1zatd5687/rY
L4UoOQ7TkIx+iK12maL08ZVFW/ZidPGGzdrv9lMe8KHb+DZ7p6AmRf4IE74RD+N0so621hjL+yV9
UKqOT0XWU0RAJXSE+Slxhml+iLbNx7YnSJDa2HDDpejhbhtXCIIU3njuqS5uWQHdbj4zAiaHFh/I
5M8Eq8+KU81yLFPcGNq1hySaZaZpYALyUhKbwouIGYdwMx50GlyRUljQe6mGUdS5RlHCwEBdlEt1
oYLemzvFYZ8KnnRQgC7yTpidnPR0Fo3FUcFC8d2labEDQMqwF+Hi9bcYf2EqjXDGHYex6CZKMt0p
irNPq4hxhG5daxhV/lhv8QLHOB5u+jIk/vL5/TgwYpB9liCXPZ7VxulIpjs2EaSrEmx9lzYeCM1u
XxRZYXkV0GhVSH/PYO3yzV1Wd1L/ZMEhU8Q/xPvt2zYvDkt2yQfhfa5bp8sscAHZh15tHro4eevj
Y9vrp+hXr2JG4PETvfiny09s66Vba1AnxB7uHdH6lKAghATpF3TeEXdcEQCEc8PqjId8JLIT/oa2
jHM8v8z9Zag4G8baomjJQBhXHgXkYMCP0wERIAgdSR+WcySFvA80bDPmr432vbH2WSH3B6L0ORHq
hw6Ou5IFDK8OuSzn6ujxvfiotCKc+gGQdf4qDQqcBDdDwDnlDoWCvHOOzZHCEYcvkBLKYn9l7P50
pvyGuMJ6G7ESMD5rvl0Pl/0kJr6SNhOasB5Seo3A1yzIgXNB/PUFTvyWJjrFVxU2tww3+CgPBHqY
QK9tjIDFXBk1Wrnw4paHxP24O5tJrN8Qo5JMtchSAXWLX99eqKcETrpANVFQRpoPi+e/lpdF3sRe
PwAeHM3ztsixDb702kDk6c+XZi3EebPIfrAtsMceDDH13xtmxabwd1PY7v/C+oZF48tn8dPiIN90
RHv96PkaVo6eFHY2UrVEF2wjB4OrFOcjYKZxw/Aen5RCNOU58iX17DXgISlr3Ix8sQEBEoeUU8TC
iWvbUjM9CX2PDreXX+9NEU7thXNNUqYKtqfA2S3P/Pa6boB6105b174NIdRq9hsUFrfhHFpXXtY7
Pf9Ka88aWqoYnwlj6whMlsdsU4IyXN/I11RWYB44hFOsofnt9m/M6oTUnNW3ZSMVLgYs6GUbi4tc
qAFksnkeAPOmVgVU6rntXYjPH33qbdNjR6vMJe5RUTrhqzMWkRyz5LrND+N6d4X99G/U6kj3yjNh
S1M5EMWBizJaeXt3k9BT2+F3Uoyl7FjD/xvLL5sphhDbK9A3IofDCgDZ+1lT7J/samA3ayFzAYUA
PIZ3kVCWdAJsgaAnQuPIvaLkBd+C4J8aDag/N7noKIiDYPQ0lYbav9Jttr8s2fGNnUHLRHH2CrW6
LUyfL7oOlE6xBe4PYvtjHT82vliTsJuBwvS1Ps4UcdERzZsZeFMLTxUK0v6eJ+5PtCYuN1vs5KSn
lSRcx1CDBbpUnvpEMTEhxYP3BI0YJNIg6eRj2Me3OcFUjBB4K85Tafmeqyv3NR0/lGIJ0+tNgwVx
/YuUeBEiseXfU8roOEtvxO1dGS6w9VN7oBH+HFU4w7rqIyjgPREQME0xS8sHSIoq3xs8UdQQkJ8l
4N7jQFTU56vVwrKEqtpQXc3sc6z103sQac1JuzlMn2uiyBVVaAduQJs7y8WfJvnuQWM3UQA8euWX
LsHuWkYlDz6Ok3+POvawXQ3KEPl6sM6Ir5VKP2S2n9QvlAw4w8NIad7omt8uNYqFhKMXK1OuVmJa
5uL2XGI0Fya0ZpthSzVnjlHUrSxxjdSP+iCogb/TmaKicPTPTB8JQxNufxgTccOiyKw10amGhgbW
zAR9ehmkKtoKLfS/0LnYirFSTqybZuQ2Nzs339ThQu8eWsRfVk6enAXhiBpJDv1h8K/66bFq5N+h
kxKgOZl2j5Vt5zbrNtFh8fXLV9K48FecshefP9HpOUzfSdqviZfe67c6n9UmT0byUQifIg7rFRLb
yzblJyB9knBFd4lVq8Ucr7nKmODUONsnA3npy47AF/ZpbVuawguvkcBGLSJO0Bgp1Z3YnsjKTF12
vzMkBIz993baIp5sv1gdEYofZYRzidK726u4H99nQ7BL9Lc0bvIibouP7KRiQi3hdQ+/31iZONbL
ZzeYRg4ka2DxKLHX1ffh1bRoIcDHzEb3IsjjlP9xAN5aoOJWt9lTrRfA7e2oUC4JfUdWMnSfU3zu
LH8gRHERRAETn7fCUIC/3JmW3EPKNcqEyT0cqIa8gwJHJn+3aYbGgEKKG8ha63d/SYrINwrZl1cY
Gu9uW1uWvx/yCj2288HypDOb+N9cttNe3saZU30F8LIYqzVUiEOW5Sy7Jlfacza9LIJgkHqfp/jn
DrU1cRMEcT5IbF5f73BpTiUk6cLHvDxeLZh5SSGT8fg5wg2l4eT4JOPSboH8F6YWDiCV7V6/a7Oe
PbeJzPUxHsPl5quMPaxjCEyAWeoKGzzRT62aTazJeycEn0MVmvnv/9c2AMfswdPORAc2pVbxzX0E
VnuhYpfJsMgVm01LzPWMaVu6S8PmWdG28z4RUvL4MPwSRfYRZXw9WenZ/PfiEufmc8vCjlx3reUv
MQSZTaa790Yuj/8Qi9Mn97jPQA246n3LDYoMN0LMDGicGR3FpQXXWdZPrFlrPPytgK2q4lan/P8y
LUDQ2lzVFVSIImoB1HyyIgFFEwjwjzMgwWJl37zQ7fOnuRyytxb3ojC7vF8Ut6cjsslErRhRphuv
vPP7jEdNPGmqKfYzMacjbsVpQQjtSwPf+9Wv/PSKY9DNqYkZ+7j94zucsPuqCpcCZ/W8B81fL7PX
sKp5APT6NL8oCfV75psciJCN7CsPCo0j+PLZQqPbbBh7MnND1W11cSrZuMbBnMDFPvcikvL5J62Q
IGLeCmuUl/TaXMbbj7l0byCfsjmzehVWh7XQilkelbxH7avMPDXzP1rQVdu0NSLL1h9tsJBOaXmy
j8bmF77CS/JyQFjfCSXJ0w9AWe9cyvHPQ1N5xxfiXtYBxcMqs0DeSuc/4GuJw8slnt4+BcK0QUi5
MItqw4SExQWaxaDjU8kAvYBFQ+lUqqngY2IfVD0WlMkdrlPfZhPHKgjROwL0s+VW1QIoOq9t4egn
zrDr6vsxCRc4FzpaMjsQQWAcGKj9s+4GABytn6PHzJNTCNg/YyqUtlHbVEavg/QloDO8HRtHjVEa
P81G0nTXZFzbUNd2ipuFYQvU50M+Eg3IahJTUpqRPCRuWlUxrf6h4W69Pz+e4XzPS4D6jJsOEOXN
gAPDq5PpXTqT6wjWYg+1gbei98T/RlXnRzdy/L3ojjbZQzhIPgeff3YKhLj2nDpdB1Ns1YQEDRpc
2GznP3xUYQy8RN0tkP5GbLJfBGwU0hOrs0O2EtHXHSXITXUAG0FhR+adqr29WxEmzMtffoqwmbAW
aBGrfpSei25UaL5ZTpFnXE7kcjDls8iu5cU1kbNYG798/SU/Io/m0zAPQvXyz8FTgBxOmiMSEAcI
+DfLvCB/nuSNWW+eOhlsoyA58hCaqQB4Z4R7nzvAVyNaHafpfQffFqymvNQf+qbTf7bKBF63d2vw
TrvPz+3Mz0A5XqMStvFpqWhtW9NcCSwAohrfzp3m+gfO/mBiS9f7v/ZuT6NR2nHFiY8X2D2gVhKI
gRb9GPFFIBXO9wPtYg+qGfdez3a7GtYjSV7DyFL4/lFJr7utt76Lp9xV256JZ9CNqq/1W2hoVDS4
Rbsy7mFZjKedh+5TcTjExgb6Li1IZ6nulhh84MbP8Nw0IR3fBRpVQgJ9ZIIUAwfv5GwAQ/hy3X/U
06yAbCnlSSS+fp85Lpnw9ol2ZAh8AoPpMs5AoqjJAZSYnVhl4tEBc3XXRIH7Dphg8hvmM40FnnR8
xqFJ/hCCEPBFeoVrZST90CWY/pzlCsYa/H2A/zJbHy3ISOXUOg7+zWrRK/IR3nSdkrkfMbRqdsX4
AFvsd5jp+iC7UVUXGD+Xxg1oqNLWTMvWWO5gL8J4+LthzhAyPtD4mYpjdady4FULvCWvevRbOEzE
o6qZQzVN1sWPeDTSTZ9OKs1F8T+OmuP3FYZwCOCSXPa+a4FArdm5jRyyvp6DNfpuj7diMb89+Aqz
uUrWN3xWxend7nWccnQeGTrtn3Ln5rmmmaA7vXrCHhCAirdP+hsgaVwP6fn2mVoZRQZ856E4vJac
kYsmGK7f2B1Tkod8FQHQxAm0STiCbiyelxdw9f6z/uxIHRrdJptY6CUxdf2UKGRZ2nyXGELewcyB
uyNtVU5sB3nVFlHyPthKNU6LM9I9JaKP/qfUprd27AsWOmd/ubu4MnvxAnYQWfD2Uga0k0lPyqXw
GuXut8huNasQfltM66leFxtXkEvE2Ktti0KFl5dl0Ag3FTcPkAHVQ4EFcRyIMVb/+o8kxLhB97RT
+mahopVydw9HIR7w1PlG1PjdNDnfA2gwytrNPC90T61NNR5ZpJkz1MPBYmVNKY/HhUw4PrR6uhLc
pJGw2N9nWrJO6k14F4j5Tc0VIA5160c+uAls14QEvVpS71Ku/t9BN2Mu/moe4mILpN91NW+WPwkW
4TabRSJo80NeBBvAKLVv7dw2GzdLLTe5NGhnrDOwN1RItouKMZxFjBNTWG5yYw5oanWX3cKCd213
Ly7SP6pTutFXYBXNcxnscDFzKZ2HvHuhZvp40/FHmukp5AGmvT3ErAxF9WqsMV1HMFUpnP92uTnZ
Zm/ozEbt0WqFxwwgmNs+mzfTEhN1Yqv2f3hx4+axL6oG+hdtmXAKJHTwTBpN+V5KljRROiFE6n8E
onzkdejzUUyCe7A9zG/bX/RqzUIWxXtV8sO+2unjRypvpF4YjbLkzvjz2kKO6qXapt4Xfdl3UxcQ
p2gp3p/lUUM5YAZN+g+GuCrA0A2TobK0AVGIAejyUDEF8gUaTboGTu31uIgrN/85bNZxMuTCzNR4
eSeZZGiDoo80WagKV1QMn3yXx3XlvaEgDUtquDbbuc5TWoZ3iyLlh4wV///eIpr6h0kGtGRd756H
uyC78FbwTvw1apiaToHKP9gv1UzL7c9DXAON48dNk6D0HUeQrv3Cuzv14H7Y4R2BWnN1OVfk10Sp
u0g7HuWnxMp6AT0bL55I0oODS1nUnN1L8qXTBDk3FPDcxpeVOPMeZc2SEUmOJQo+XFJxzpKF3JlJ
xPWq6BICjZv4iwbzYoGmkNXBoV5+apfBoVOZz6tO98pMHbTykTBShXR7HQbzj6RfqDEE2sYv/YM9
3+GsK/mYWFx9nDM/RP7LEfd8ntVWRzklhlt2V1QCVOPFJqherR+ImeLa06iI0d/kzdKx4q+f2FML
BCBFvNZJttTlU4LFX0ic2LbWbOO6XHB4rSCbWwRNsqds2HCiqSlSl/zFna2z2NboYFAK4g7JK1BR
MnjXX9RzJIrTSPlQF+kXa54kOAPq+GQ20qY2RUUlz9cY820U3NcQroUWBIw/n8lKyKVGg7Bh569E
3qW/dONbH7/sNrDgWG89fPCFtwOc6tUs1Pav1D2jOC5Md5Gjef8weM5FKMKMcllHAnPa+5lOItvL
7QBQp3Srdw/Ga1QCtLMxuueMZwHLQRnLiiGPPYA0aDWkH2iAt3czAlVkX+GjySMBf6o7PXUbapoT
/oKfmltC00Dut+DOZjRRIvp5A7YeV46f2vX28/GRbPOWSnMzzmDvPEYZ90WeKoZWW7v1kTE/GeDJ
vI1lRBupP6VpcbuZsiD18Y9PhADLZrBS7cG2Vd3hpjqriwaxdjWjltm1IftJnqeBqyZF27MRzO+x
mNM7V5+GCnX6Emtf9vI9IBWM/os3ROajAAciTpQpmQkiiDxqmS6E/cf4VpkQQdH3x7ycYgWWAjil
cbWt74dnurkG6nqBrQtF0GxdIk35slVAfRSMYUeWnJHgKE+cFA2wRVgweZwqBL8cZZ78/d8a/bdP
gl/9CFhVTNjMLnGhze5UC5U4JUGUosnhQJ3Y3fWwak30Z5EwqKsFV81Wj6DdJ1nDyqcxolEO1E4d
0w++/xeVHdEivWyu0mLWerlmcxzltsR9Ua32tWXYjquR7GKIVBjXHIBb2co8KCF7M6c1n2vE4FEV
Foo3NsDtTISfLYXiey4rwcnHtI1E5U7r4fMqQreD0FmHvpwqHRHOdiJtFZt38ScXYRRVcITzzko5
kyKX6B0txfb+1qMt9r+M8MnRqGrej5LUNn2ZlzOoLFtcSJ4xLsxXkUZvRVu5qw4N5ibteC9jzWIt
JIzsu7YWi9QQgkhfcZiA4mWswpqtx3m6aGlElvT3BJRfmt4c0CsSyJzbOYl5Nqlojl3yby4+2Bhx
1Uvcn4Eg7FFxt3oZRONjJ/F4Fn1P48AhXsxxmqWQZc54Yes+f008Bf0j1GxLuZmV+XwW6u/tDQjI
E9BPoaBoYop4JeLhbjkrDTW4+Ci2Zp13EZU6BaeCv+YDs+D0cZptn4W3I63mLTE6Ll4h0wPW0Azc
Xoaj/3domWUJQxYwk6cqa4oAamSEUVRzeblG0auZKB/OpXnQiDICXzsJh164cVb8I9kOAPwjg5vL
hAya2W2NiazJpnSkRdBg9RzhLwWk2+W4i2/NWeOQN54LEp7FAqPSWPnOFHu7WHJzRhSSuejSGQRy
Gd/3jYYBx5tKCNOqfJHeYpJU1ehOYduWDgBKp91JGL/RbcWFRNs+5VBq+8LrmST+MPpDhsGuAFeT
afr79e38dU1SKD8CWxsqh3Eb4CZjfMesWyY60epyFOMARMW/GIpCJyGqULU5P4rr1RDmn4aFBneQ
5LHI+IFQMRjceTfKZOngJda5xDdoVERfWgMZf1umeHECF5/ArlZi/Ghciuhrd0cGJw7fkmkC9Vyr
jOOJydC7hE6cfsfD2lPiUXOQGPnLTIzysZ5Lmx1IW1uIGdNi4vqXgUaTpD31yO37u6RS+edRBdFy
MuyfEPV+vR8DLd+BNVlORhBMlIuAan0+fiWLI7C+CpEwGsJLpiZ3G1lD7MVHueXp2y1Yt7bWjt6t
3RuO/cJveEUW64J8h8YfRWk9mUHtscDHwZYKqASr76kFuFQNKDikEZp4jissKl6nRsatMDelJkg9
UIlIfyXxFSd5gVNqLPh+iMDH7YT+GMMr8hZW3dkhAUpHxvjnJy4Pu+cIRb5pOfGqbtzl/WJKrqNx
m65i7FZUVKu4WQ0oYJl9q9cpfsDUZNZSNos62YRN2HcpV14s+FRUaOK+4YDOaNlrnkyr3Foq6MzD
4ZDmum4eP2xnT4T0NiiOR7Xb2YYjtau/y9TIgAY7wDaCqTVtK50l67e39hTgujM4USo8sz36bmjP
VtJGakmOU7Q61SD29ifKIygB4f3bsVrfhu04/jETqg/YvyNGsQTedncUjn1clG9kBkUnoJ3a1lqj
axzNAKxTKzhEjFToD1dWhHLpoTehpc477wbGQag8mDNkpmLX6sIa+JlGTPW7tUg+Q0m+Y1F/XmbL
KJXJfYZ0gYdmJgpZnf2vhI1jhsqh1cpydGH46RpHwrpFeDw5AybNchMkN18biL9qaKCtaYSrkgNL
sm/PMgj5hl6N9l3g/VPVJMy+rar+tVB6ZY9bYRnGIHSAkhJsH2x5pFOoJtvPC3IlKPNktJWR9QYz
BLzhQEWJzuUCbwCDMy/RoYqlmYcE6V7XhNBoYoftaiIW9kBtMYMiBdV2qXsSpiq6q+3zmD4OCkpN
0gnrsIotmGZUY7AfTBUnHlhJcIbuFVlIxY3uiaEsrlHbSvyDfJo2MaGwLKiy5FSAnrztRKLWkxjZ
LPAsq/ieGWlaZD+yUMRZ3e7z5vZ3Ewkq8MyKR63kZg5duToa5MO8y5P93OusgeMZr5yHEyg45UtD
eSR/fJ/UF9neENPQyosVCuEGPc6a+vmPK7KpWPiNCCFmSTD5wz0W5Sk46YrrQSg7T38E376fOYSI
9/oVasIPANbedW8Cq984wI2ClbE7nirsnD2u7030UYkLFS2AD/VjHQAOFqRTllhsFhkPBHe46Qx7
Gdzb6BeO1T+mbg3FqD3El5pfwVI82aobbUQgi6WUEzkj/0S7XbrHF0qIwVP9vYOJ2ODMfw2puGY4
FrD6lNufw2UllJsyJzMB/5BO55Ip76TYmUSzP+jZrL0Au4WjMNX4VKKl9YWS9BJNHfzzKWhxpBGV
IX7W8HWE8i7st80LfO1O4wyddaro0t+LmW3aEQWf7xXxP4gcrmjHFoOx1LHhP52b+2WYgr6B+UlR
709zztWU/jW0u35h/P5NI1dbEhJsyKcZboSVfhEeacla5KZuV45takxCoY8uOCO82lIzwrxIkgpr
KqmETfx62YoM5mGhJ7LyrPv40Z7Ea/TTZza9GuVJQmZbsO4QP/qZYWe223YiBrBWe3evXuP4GMHB
/pMj3ey/FzqzpM9lHIqE0UXTz9u43JBwNB4zBesTkyvd6MusPRBbb0R7p4x2s97qdMl3l6sP9hEo
9K13V4UoFrH5RoBFbeWnGKjE/HrPtv0Tjlwc4+7pHqrPzTtiZ9/tTbfXLqsB001qv7EFWWBlff3B
Kxx9+1Uf2USybXp0ymIu2cB2X0LZnE6vdcSyH+9zpJVchrEon09HT356u1JOanE5fR9BD+0xUSAA
j0kVrjOH4MMEDgeJRV6WTNEsu71UA9Ai3L5v1LSZat2OTQewVvfoeIWkdeXMdo/pptCG2np4Bt7k
zbYusRhbmZUu6sD8lso9259Xa3DU81yTPRLVQY9oHMrGcqFEwMi3HGgtKfQiR3ITPNzQn/ehmb0N
ZqFHRlLA9DLsufPfj+O5dCDju1+q06Ubeea7JTTX5qjFXoecNagI7dcKjMnCyVBPfrYofs9DU5VY
STWXkvbFRgCBkHj4uKeUY3YXbbvXxSQOfcDKVcmBA6x2lYHCHpo6/T7LYZjQCdG4MkUM0HoLqBpi
l96mpXhI+gfpjT2UHxwoEMCJhdz+lc4TRLMzyVPZJ3F43Lu+3xiN5mVdkt3c3yCRp5q80XjUgUEL
E3N6xFLBB3nIb7m4wAph3mom45CQsInilFmuflnS9VzTm6gqEAb5+4iuqb9RxlN0WXdf5ig1NqCh
ZEHzU4CE1nQItg2/LpbvGnUzRcEMQTtHjPX9PgMB5A1aIdD6yVkQbQO83ZtvPjBXG4rhumIGsGZo
KcVUnFjuXgEBSQi5Bi0HNu2TI3Q1+lBOb7xQmcgV3rLTEHx5EnDyiuybT7D6qs7pmf5+Hrzj2oPr
LVuVC+4vgGpyyFw6v31tVGNC2hiatVgEtXYVbEgaWZbQT1EMwyI6R/S7rYMaSaUDAz3gZrOxEo6X
VKGseC1sL1fl63VfMICCu9IjhNGaZHGyTRhBlTzjNFF0bxzYwBKexUrf/eVYnInndWNotBGGA6dH
Iek/weX/QDpezdOqosmNlWQsCwfcn0mzpwB+PYASZEmr4rEJbimsMr6mT4/EDCyw0mtbeAbUZdf/
9m7zq6J19ANeXSKb9oyBBl1kygb3eRZkZdHqzQ///vK0Sjt/u8PB59dSP7C/CD+FdwRms8DojH9y
rWA2Cb+2ZKwpPx3es6W3SIVHqOYDihBI4M9qRjBDBK7E6MPJq3HxcwxM/P7MrDC9mqSgO21r3zLP
LJy0JNZB6tANA7cINiCoLgRs4+CnKuCS2ASpA7Xd+BEvjMeKjZmvxmOkpiQAj0jEQPZqB7Ihpg/r
M+gg57IA0KM6XFlfcK/Db2+F6dl6DfbEtZ5FIs8bslJnl3XTeDEfmIXLQIpET3HbZlSAxrFxRwyy
V2nTxExAHbg8PV7pS7t5xNXDjOsGdfO6QLVSlxHcpnt12mM80d8HW28a3DxSalzlRtgq8fAyubMu
KfxLhJDTip/k8zC7va2RnzgBbCc/+V+nrrGvfmlUvgpaIwc+vxRv2xzdNLAZ+dq3+EUs2s7wgLpg
xOZSc4Ur2WcfMXCfKyH6A1qDUNt4f7Ch5SJCbiTEA+4lWoFAstQQoB+cSogMW6FsViJe8yrVFYcX
d3AtBBNTdnZznXrryDKApwy+v9ZEx5J2X/+PxAzza2D677UoiXanTamxgj0nInHYYCH/bk6qeFw/
ZWpHr7wTICLWJDgyohyw/EH4ae2i9Mq96EYiJyLysli/UyRc17SmmU7SNJf2nYzQ4pb4w52aYoiC
WtH0Rs6R1vJp+JvIiy8PobkOCDA0KpAz3wuzD7OCDKgF4maQt+DMWmHz+SRYtdr3+unOFaA/PoOw
fmOVvHo/AVoced0HPNloPdRWtQ9jGKdQdqbfCZb7ASfdbsOdqVhH9IYR16J6R9CGdUX8hYnWCth8
qyecwiNEAGNGOEmgibKGco7hiUQUuE7BXc+baghfBf1RAZWxKJ0+NmuEvvbBdylFVsOc5Rqqi3IV
C4EiYGt6NVbyPCNf6N+Bx6PYmTWD3gO24h29kRbSDmhRopk1BN6jMKkbbgTYn0k/x3dOcAihc9Py
Uv0LP8yNfYgMYLylEvpRaJNdd13PhpzrPFvUlM9/GVq23SyujLOA+9P8VRVjuSCOQpjCTWs/cBi7
oAlD29tVqFq8NRGqWqjlIzGuHVsxCtVusxRZjG/qw7T1fCa+bFxMHQ40I3x1uq6qGqYODcDA6m3M
ikRB4oCV4rZcjm8Op3Z6xvPpL1hvP/vZBr4k8L/iJANTAqOrUIzCd0JdxfDrr5vSEauIiz0YtlrL
tpbLIez3X4uCcJCN5ASfiQEA8atd5z9TM1jHskt2mBBAQw/FinjH9bRHtuu2w2k28X0sEWpJ7WU7
9xRa+fBMqUozaCiRvodymECFPLWxZiOrXAS6RRJD6+XvOk8GY0TraqiFdoza58KF38eBCJF+22F3
u/BH82uXN31ZtKXvN81U2RlYOpP8oxxduRWoao85l31b4llBXqhnuOHT3tywbtUTiA0PKIzBhBPs
PMP1cR+DcJCeB2ToyIzpG4bm5zdXnRpUyofDLnyGtwEMxWBw2gWawzfyc03842IvCyy9ZBplSU5x
buWDMzIhwXGpf+RmmHJ+G8yFCt45DZRHpBGdZCl+l9N/ejAR7t8/jOehHb6Kp8Qs+oljo1gAojKO
g8doZZ5pD5K+YyEtkJcuoeNxGD5vwk0q7eOygYwmmIw6DfVpdGJ5XZUApql6ep8jZEzJ9uUNUPwD
Mi0K4ygX17QfyAvIlQNs+1VGaHjiBaNQoyXY/C2JmVtkiXWP/+3fzPoNNUhrbhC8jO0Pp1MMhkuy
KRPbs3vLYLqeXhkecPJFTn1uuOEl/AXUICTDBH2f5zEoDl90+KF5AU5Qll63B1yOzLZEa+Jhdlpe
0Dwu+2uRS6v+bTkBFrE+GgV2qFKe8EmetH4FUYJ3+5ySR9vCZI6/SvYlgL8vzK+QCiq9F5lmuE1N
aBi2jNJ2G09K1JztR92Fb5vTDrFUrxljK6/et4iUcGJT6voNrMGWhN6HhVhRB8mpWxq0jTAI8gBH
3WmogH/YeJrOVGM8kAWEzMv8Rulw7XBaWKB8AaPusRVZ7e0GB/7tVQiGYQ6y5UIYPTWM/142Ozvm
aE0gMtVeSkKJ3UlHnRvDrvUDAcLSaJ/wMopnp+Ki49riJ1VIZhr1pcnUWXtebOkE1ZBrzuF/fQlA
4V5gik5nClkNeG1MWmmcOfXD4GMMffPglQT5kGgZMevzFtadXjl0z1x9Va47SP6AiXZiBg91nkmr
70RXjzic3+3PlrftGSGh8xbm0S2vBHIbFQkaQ6ideFZ0IX+Pt13HIrMinCx6P4iJ4177wstvQdLw
2PvYCsSXsLQs/o2j+mR+vzWGmj2RgRAycyKb2RslVEg52MKFtaLbkiMc90PEtHqPDgRpSaJzPTER
A3g2DBkhDKTddtCtF6R10gA2uCuil/5Sy37PdxqGmYzvylwPYi9Iuu4sxy1n7ONRWQFmsUddrNXY
Waj/t9ChUF2YbcRzByPU8TTtZXqWYv5Ami7ycuG3KJUZ6qdMjkGsVvnzd6F+66Qkdg4bENu6XUAp
CHj4fv3lP9di2NUfB6sO8xxEhAzkUHahe5CbqDZy5g1Qol47dK3K2gjXFtHtW3AJTX7SnwBFTnWe
uN21b3qGTntBgzDMM7U/JtDssWly6K4U63qkL74tzVnpLov8xGrWjNTthQccuW3YggTVB2in/5SQ
jh69L3sR+NTIHjXaTfw3/Kk6mXRCAhUJYR3jMxOwwwvEFrs09qGq2hJH/TU3t/+F9xfm+ohngsOr
vYed8HKv12OHIYxlmbSIQwOwc+If+6sYjQ4jp4UXud9O8FXHP0/E6ac6KuqRki/Rxk5VQL/frvzz
WkfMnRev3hhluRRlvDIyYYYiFWebqrnkgNwY1tSKiTfPgLxUqG2RDXyoKuCVM/QzaCrv6xkB8rog
Mr+76Yj4IkrKNWkclCfjQwWPtDA9r+iNzn3dvdInvlr775mqe//k8KU8bN1pbfsd5O/8nB9rU59U
dZz3CfIy0++rIv8aacb0ZWmCRS5xivnaWOVA/oL4fiKUyNrrLCZDHOHzeKokeTXxxP7Q3NE/RkwJ
d4aSfo/Tl3Mlt3B4jiBI+8J7P1tU2CfVeMmyu8uammb38l34eQ8dQoCTrhP56JZrtfRTXEYFc43H
M5A8ShIFYsl1aKGs/fjgo8Lx0AKGXrQYXPxi++xF7ajnTWA67RJNgTFjLLnm2LoC2+uVerJ6eR5J
TNk2jJ2bBQDHSmdO8aLFHF8HNvSqo6WgE9PfqEiqFAqnVe90jo6o5/bPdShb7lrvOwICTHoTdHD3
cSt4w0y2igT8OfrjRUCJQ2JNTel7qLjCFhkv76j33iYPnYgNEXdgI+omSRND4aAIrutthEkEaTWG
cHEKsKQUiQl7q9Xi+0Pv+3sbOE2XQ8S+6N1Rb1oz2yOV1UssemKmRCwUqoT2lp2lGLDFF9gVxM+4
5Dr4UR72GcFexKyevs0ZXumT99/R1p6gu1FaofjuLD5+sh1f+FjxxuCoxdpO5yKE3vMQnu6ZL4oO
Vmf/j/NUrV3vZKIfZh/CUzTSToQyaEVo+X7022xzXVJ/HK+gjeqfjWuS54209d/uw4cDuuywOcCx
e/5OYW6hNqX1WGbJXXKI7QkzP5pyzlcddEpb0bzkkYI1YvjcDWhC1HxUg7EWDbVykyaMSX41yEYU
375yQGiiDeWQI4g5WIqsS6Oln0dXAuhHNN2RfRjvWaW3tVW+7WN0/OmDBeAVI6eMwxWU3qmOyY8U
ADtBUbY9hk8CrBXrH6NeDzs3VWzTmxq/1Ihv/+UvbktesV8irBySVHvTXqCGL3qK9H0YZNJvWrVL
D42xpZ+DBVke4W3ep1ussmn+mhXrHd7l7vF67hzE1fwr2Llw2b6lsAhxznVLd61B5q7Er5HiVrGA
0RuG3jDNC4jxuxl8FDsHX9SYOP0VoitFnPh4dipPEAOIPcs7nXswn7uaoyNzIB6rORDSAXPWT2O5
hjnCrYqETnGHQOYF6V4Iqe/qJdVQp3Wf2NJuniurEY/CEwqJzwCK0dBMgt06LsQ4EM+inwgfjG+N
OZWRG8Y5lAz0mSjgjFLkhOtaFyOQrrdFvCksEN4MgKOLdMC3E+dLtBztkMiuGjC+MenEQN45lBE8
6+2FV4929ICVMNrkrYDf72Eu3MuqXS80HVmJMv0HUyPpIk7V+hyMnpdOlngBA42zY7xhTuIu+BoE
zL7BHWrcE/m3YK2zJkk90AwBe6otYArMbULljhkbkNBMWRUS1d4OPZOylwCAcKmEroz4nbWdJGkq
olAszAbVXKUQX4hbX82EXlGWtXYpuVS7p5GrbRPmp1X+bWw4XCSj4DXwMb4IMg+KbWciQhv744I1
1s8lWPNFNKseshJ0jIGtxd5hJAwMy1ej47qQWNrQTQHBYE2Sofdu97xN0oFQDT2WqDPGRFBgqud1
OzmEdIEQM6/ZGvRxsHL8QZEQhpeU+voMnEOaa1DWXaMuUNPAHKXfL5USYCBSP+uQaKSYjOAKsx/t
vkBzGeZ97usiR8cbfvRWQXrC5N+Uzy4j7Pj2yyqqHTZtj8i4yqcCmW70qlN/Aq5Ih3X1nutGQv3A
4kxjoVES9Sb4VuMtdie/yGqBgvaGPwi9tL5Q5H3Ls/3DaVe97GE90lUbbXYnhIIw7JKIL+C2U7A3
RRCIqxsy/24mZW7nwY1AA693TaV4l4NsD3SYt5+nIp8ouQ9PdEEalTqVvdcHFeOl/tfuRPrC+ZjW
kmnIlFgDV8w8WIKoX9/JVPSTvD9A5PuuKTFj7JJUMc3RRhr2fQgrJKd90XOhNwNyb/SJcMA3tZNd
YDgRsCFnR4QSRVRFUMSgVafWtnTsPj9qyEdbmNyVQYPiQzoUH2kAUM5WIGaepbX7t1aLJ/zEfozS
49fz6sjfeu8gEfXajb/3DkQc4jeoaGyNTC+lm+f3V+bLvvDxbAJd1sv1hfkZigIksKKV0nQMh4JK
NF+S8Vf3o3YCFG9syhubIjlEKe/ryO3gjx9i6nqss/RUW8zWIkp1TIEI/kuu5+9OIZXnukVQxR87
iqs0oFeUXl6Gu2kVjvEVDjO+4tarUK3f1bie0ma6eYHmlPM3D8zEHYAnuqVc6+Uvlqve4ScFinG9
6F8C6nXkGeVid8CaiYKPbhbZuhwP+Q0OpEoArmpofyYkv9SE39lpBcRy6MFcdBI8cBDJcKwGf2eT
zDKXISQ5f3V9yPwhQQc0c8kTryyzYD7H6rvW3GJjk1LTsQORS9qMBXUpe1mzP+CGWYbQLuwrj+Fq
qrnkXC6iydh3lkTnHKx2GoVAqoF7Sc2yfNyQoJ7c3soWkK5rMqtloTuatSHXlcNWtf8Mli5DfOZx
H/rT1fifO9eZh2o9KNY797ugren0TxJHLalf+jgISqq+aPU1XkjwGuzYpMztzjD9dfUHNvTPe5xd
fCic4ZLeTTnVPYGgDMzG2Wi6Y5NxgYrSqzgRDyvAExRxRrPksZLNGsWX7guF+J/7mQeJnCIhH0sZ
5rLA7ZH9TX3Jq/z0RFnD6KKz3a2Gu1X9KY3aIsM1AFySUXcurn4uDxxxMT+FWa2ZtdkySIzfSgzh
taIgd5aIfS7c22+/V5QeXDwbqBGpfT0aqgJXsNuBZKRliwJi+jg14moIz09/tKs4ws0beJyS/1tk
zZwkTWJa3Zp6hX2KNIDLOQh2drbzF1vvh/Cac47DTwsALeWyF3d2NswFrJJwbZIZ6Gc6WRQeoOVD
urCTSrMF9BLBVH8ljCWFCZEQOKvsNGdNMnVXyFa0NogOuOC/G5FMIsRnbZ5KqMcidz79PNTdsnff
/Hhqj2zN/sAu6q7Z3mS7+MVSU1HSvxhVB8uJrPGTp+9ruX/8F4LqrAHffL1oDQg1YZk7EfEoyR7k
QPR1eKvxD2s4iqBTphzjIyZKy723ngbpk1iZ2wJKN9B7zHWhn5AL6mbe5AXVP/HFezvyAhWPUXtm
YT6FrRckLDrzQHNp4z1Ags3wWDuiCdKN637qjCPArpc5ZWAEY+KveSmYXYGfs9KwTIE6gkcotITN
PLnBGJMXrI3lrNQ0vuNbcwxe88oxT/Eg1ovzVqA7ep+sbJkzwL87r8ct8PpIoAd4yB6HjKZ6jBF+
j2Ewzf/XWErCaL3AFtErLyH//VYS5SAfNj98OyGnK8r9r+iABF+KA9w4ZGdtq+85JpCRcwYlRwI9
Dy6TJmd56w2hN62ZPwdUvvm26ekZ+s/Y+D/l1hnUfRpGTNEI6o5nLObDLrAd0f7I7xB2o7gK3+WL
KNQLePvjjEeu1fCEU/07mEKcPRGKw+qPln2PgqX1eagxbyM7k6wPScYsCtzoNYBabN3Adroun3dB
m0HWca5+DEOnq7njXtEbjTWgXBnXVA/s0lF+4TkYsg4cz4+N9PfrTLw/j/RvXjnwZocFD9A2EicY
Z2Pg71yRoZtVGDypTHMQPmyQIviEkXEUzDpKNO+vNJJQJM/Kje2of2FQiX1m4wjbAWwiBII9lxgZ
HGK8SBX827HtQ38QTDd6EWwgXRJYtgWLgPKBaXqrX6AIxiZh+uVs1Ki+PvCdpvbkVJtqYwxCG4d7
BsDAp8p2PbUFUWA0pAx/tnnozfofdLRLfys7VvfJresmNyKgWBcj6wqkr2kf28Z7mOnH8PkIanaS
OOGXBfRWm+kyARd99GjRQTIRRYwHac1mz0V0OtNfciJeJTsRzI1gaSNUtFmgMC1T4Pc05155OwbY
IXMPmwRQOg79gP6IISsJPg1uVgDEVEe9JRBfEFNIRcT/bSgeSLdO2/LQwKvGKR3+js6Qr3duSlix
vA1a7KpXQIPz4nHPd1Sft0IpLDOQIJnFHf6II1VsWCXy1yEJnHY/4bC3K7Q80EkKWJnRuP+/UbeV
2VDlHB4p/ST3zsAbIPgqiZBboNma14Ijjjsq3S9zm+h6syAPgVF90aXxNkDcOpmbdBoYgWx5FzOv
NsgFA53GDwK8s+Zk+NLmYGRmKtsvLu1yyyeeXlgIBQG96loqokKVUeZHUdjS8KHneWXnyGxAFim7
pkesPI60GQUd2mRqGjCG1ManXgWL2y2dnhcqLi9W9zjXRNrpTRCffExhcwr5cO83jKfSJc998yaZ
lU276R77554yQmJr7gnPWGqo9VcWM38d2SsH1WpsPNaTu8iOo2oyjFjzYK7x9AkD05xgdhTSKOez
kWfDlBk/J+puP0BZT3OTLrk/1UmBOpIoEUbsT9ZgP1TeKkrSUxrGRzcqy7zT549Oi/jCzcpIbrXu
iEMMUgjI3yD7umKx9QYVAxKLArwZdHgHMcyPwRylXBaPcvTeAMqc1L4nBf48g1ggxCloxt61z6Lf
gAgM62u1p7NwCxA+EAVdB2XSR7RPFNaqtd9t1cauEF8LtoWi/AUhriv99O+X9sq/WcgisoWanCp7
IRvilyN4AZlKZOaDKQHJyddh0ytDLEUmwRCLExXYrRL/JmvnvqSFWYoqqR3ycisDoqZCi3v2WMhj
HCt4LM78JhnQaErKog7cfWGNuuoiuKSV9kYv402g+IO/uTpsEXrxmnfV3p8hNgme2TahI92srQG3
CFfJZE2vQBmezNPP0Mn7ePQZg0/ri75A2nwOP1x8984W1MI70MoPAF77rTCaUo5Jp4aSLtc8RQGV
yPOZvcn9/uLE94y8mYyfDE1h5a38YfELM/+8JV+Si2p78ZPwlf0Vj4ViI0o+buPzDgxbL6woH63p
UdcwjCgNccom7zi2YAd7NhLvlZ0MN2Gm8X3nb8TmtosW26+4tVumX2Cpoiv+WxPuYmCAySTwDrhQ
yvCvEqkIA5g+3lUnAjR2ScqdD77VIsP2qP5hjrQnHpraOHkVnqhsqbuy2rnd5Ii/txNeLnHFJgnw
O+O0FZwdRDgY9oXm9c7Ot1mzaZWZhCb6M7L151WcZMV8Q2cfsxtTavba/JAHgg9cZZRLBevprV8U
tFY+/O0uFE4avZaEJbVwnYja4aI8Igxp0qqHyRjGwCVqa0rkR7IH/U+7eelav21CZLJv7nhi3Y5K
2dSRBSCF3IP0KG8Id7GO19G3EIR39v3QlIW9ja0IXLWoz9OdlAdjuojWOa5rdV753tmC8LYP87FD
7b5WbdBW+7eDyHgUJYv1fqnTpD7Pw6lq5V0bDtGEMj/R2O1RF58olF4Ccy4kHDmgiXLdYw/yeE7C
VkPlqEKcIRx8qMsOTYpyYEjwQ79amzIxfdLxfto15MqFQaBvkeEZZYleCRuKxjp3kspo9wG2x6Qf
AFXPZAeWJlB2PHV2SOVU9bzGLAtAKBySYvFdWPTtJw6oei8MqQk166O5Uz7xn2bR1kQ/a15y1LpH
7BoprWnSiHVhUJPpfgmMmFCghkFJxv7seqklYnjWgeKrZUktPXkTSB6lpkrrB7KnzX3NjR090Cq8
/mO6g8LGfmVXfj26iD34Kkk6dFw+YIcF2xB94xJ0Ik4bbzqGQea8riJLYIFcDDdnBTsrG2lp4p+Q
8m2+f7dc4MgWgCQzL8MtsYLy4WE5ab+J930SjtHUDhN5v3nyt56/8Niu2DM2Gfm9CnnX4lth0GNH
yNLpV4AqqxInAhP3UlbXZL35+rgGu0zjNFGbnvsVApVtjvfHU2jUgeUg9irAyoo4aV762xQqHX1P
7E1WOXdqu6DdBbr0Uo668sNfQKL+cLB+o9eFiEBD2OkbYWcXfiX8LU5ASEV1vueNDfS/vwGNyfEh
VvGiFImElRAYAzEBT3Z8/h7UgJN/ZNIceUwsiECMomci7D1PKh+L7uK1n3TaRFuKIOJGy80HpH1E
+RNNmgsk0KahWvTDbb02DbB2TOvzyYSLiE+UWLrip31q0fFMLYqk+xARcMsUNP97wziOIIvy35IW
WNxGYTtz4CbRBdeoCXlxTIOepXi2aqAvQ15ZMON9UQNOT1GsOD5aX+P47AfOQJnp+g53wtv+UURS
u+j9AaGUyuHKsF3TJJRqP7Uk84tw+N5sPTa4qbaQMMVVepKUXXtRiUTxSywtI1g4lTiprcXHFled
TZf+z6UDJRx+0Do/r8LKQBV47u4iGgPVROAZppMclh7WpBAyvfEUNdumxOJUsTKP90E86T0Ja5nS
HKQSAj2X40E4oCerzwAFHHHRLgA7eHH73VIm3k+2Zh0FGzttPeD/+WPzwcvJsOJVHs2Fd6ynCScQ
EeblynxKmXnV+X40P2cuChHU+izsamWM64JR3fsWwazTowPIuDYtFGlpkf62MIZ7V2Ogn4w9oIPq
hFpBCYZ8Axsvje7pfU160NFQczY3/nuLY1gFjn7zUez+Yssp1FnrbexiL+YO5Q9rZaXSrgYXNHbm
yTK6WhfQEXk7Ftkw0RH2itTkh/4a18xm68HEOFkEb51/yTY5/k+5BQ4Rk7ta+5qIDI9nm1j+VfMq
ZtW56ZeAGwqWJYma2IWI86FJ4LX2VkCaGYEa1RUmuiT73FOZmD2jlFYPedlrcCIa5kygEb+spUxi
W9CdegEQsI1NpNPMEPSdrqnZRaS3J8ajpZd6NBF4ZhV3RFhEdriQw9jPIz0+oEW50CaTwQfSXTua
KmuEs8xltscdQIFONYhTkynq1X3gLA/qm4EwqHDcWzxf6eXHO8UdSPtyzwJKt8rU89qieMybPmdx
w2Qxytg2fX6oRtxB17a/s5oZ7goy5znCgsVGTVwQlK2CacbEqk4HHqhBbFKEZk/2EkKVFajCy1/J
+BzcuId9U4YdB947Uhxai74RK+SkTxga0+3B6g4XwKkvdVl/rPEqFuvHT32cREfWln7dus0DM9+S
+1hs1GFL+nv2lx1Su1Npy9JODYoAa3sbVTKdugwRznA3YFd5jval8UbLRRCYmtSDhpvhCy5zTNS7
Drtf+6u7SvQbpyUNznZLm2SEOJZg+A0B6KZs4uXXA9ig2yxA0842BbXSBXYOrm+9D/6WwgtRvJtn
RaxysmAyY+2zBP3Mf/pRVUCuyP/rrGALA2UhMRYsaGlmcKq/DZ7Z05/y7l8WqM0dgUE4YdfrvAHE
gfIcqN3fXXoy4rpNYHPVyZzcuXl+xu/1ec0ew33HyrWhRFarP1rvlWKnfw/FeQ6ZzH1fd5REY2lS
k+GZuZFhTuqxGcSxlC0HzZvLDo4e3BAGBjo0JJ0TqzdTBBGTnPmaUW4GTOtxzZcBEv4QlUQ2TitW
DMN2QxoB+aK8htiqir07uYkaetnhXaiqKOBA0habrJt4tGno95p8YPJwJCRfJjMLTleXgOBSZSbF
zDFzySsm4ooR+WCWJ9Jmqx4h74jn6DzIuPcfM31qKL4WCpnccf1HqRdsntDXXgO23PxCH9dgOvLu
amvrN7uohsElfxzHF0UGK4m2q96upPLa3vkgBOjeWQl7tVQrOq8tQMa/IHKNLtNOlSzgF6s0ktFL
duiYHSNqewEJ44LE6WJMHl12UYfbdohfU/2cE/gCioGylnEmE6CCY3R1FzrZfbbssuXo/g1fOGb/
+1Rn3jUlItoZnGyk1pafersj9j56Nz7q7DjzhHPGcWviiawOWW1iYRT3a7jnM9Sy3sgYPl0UER5u
1rE/giFtqIO6QMKolhuswGqn5EtdoIyX36rdjlY8XoMJkyZYjHB+9s2R2H4x83oCuQzc5guVZ1HI
9oix9MM4wk4DtNuypVSSfPB+hDETzwg9zgi257ldlzT9pb1l7bGV8vs6QjTW+r+HN+xACNVs5/y2
VXMA7bxx8YTeA331YmE84EVHiGr4Eq1KmfMKFfPAs3U9MyFwZOUoJn6l9iQ/llmvBpbkTa6lsXwf
lCnphhUDqDIlqjKx4Vdb/RroK7VxTXOc45dw9TkG5qtce0pu51oRS7Y3xTFUA5I6GkalhsECGHEm
Ji+3zbFOyw+S1JjI1FDJj9u8IFXMaggBl8gRL7r80iyVmk3gkctN4rTPA29AtUTyGAQYYyIbZMp7
sijgCESWv8umNR/xwt4ZzzSdHTQgQeOQHWBVspigzDgUuxlrRLmLE8icQqrrmv4n2egcXyOC/Y4z
4n7ag9qDD4BWAafi1JBLV/96vcxzfMkDNdCdrt+S/qKmWTi23jd9AOmxMr0AJfn9hlrG9XzDf15c
cXgYgSFFXwbm4nt/xXI1qjoHJQ7749wQ77Fqfn/uYWcwbEXtotxiQUKyeLZA3l4Mu3skPpQ3HXD4
gk4rtZygTjAJb2BGxlKHrNnGDjIWAHirvss/yMADuuV0oIwIP1IvWHBIfr+CdlIEOu+KIs2EQf/g
1Q/YraomIdldorc7CrbNGfuClzr+B6JQcS0Zmifk4wV6q8v1Qa8ly4ruLzCm4VbrCPTt+Wh6YzIV
i1aNbtJ0qYzRHHugptGg1DTut9MR0Tq94tKWvy3x1MICBEZjy+bSjgXePt3/9kMsfkxJBhSDzTO6
xqwt3O3EkuS4YJ+ixfPka/zwN/vL9weDt5GAVRROYkZb++SElDpHmf1PEvxUG/2neR6utgAIoaXG
WKA6MwajlBBJL1FkdsS3eyg3vtJ/tEZ3vyYu3fNZOa1bLi0LDGFKdYML84iSzXt//tSoc3Pcp5S7
Y5SVxDpvIdo2FdqeLrQ8OukjE9n57tysANqrtgEYMKBwH3u3HXmyYS972LtfYWtJzxSRQYXQwun1
hCrXpupL3Tu8/7pMB2IH15LqsGRhT6tHk3RmYHy4ckqfhHaJ+0Z11xN1ZGMcq03IJi3K/hiTR9Qm
SyvDWTqiHJQK05p9gEuu2LLHEIYivX2YKj/YINo2oEzfgnKhzCJTmub8XzHzAkTEQG8PGzPhOU/Q
ePblrjyrXKaf3QynHkWi1RGOBeIbh81p2WPUHNLCyC6OjhHLNBniIecYJMT1dQ81IUmuWa59HrCG
wJAinZes2pckNjLZ0tJf40TtUytYDDD0M4Q97TZHIVHJZWc0Okgssaw/hX0S83w+KSBmjXyspA4T
AMh3MGpMwWIcY37YBuCNz2p+ODY0SS0r+FPYdDgDtKQ1BZgdCyd+mjGfwTUTSFTs4/QThwX3haa5
MixG47W7+HJ/FuM1oE1CrEQZJVaZS/JE1B/OZLnmQHCkxn82CNlvs97MLgpTnRm8NS/2XxzMSj6b
TqNq3189uazmS/W+FSgNLB4gqAVIDSPe1qnF9mS8hmGSfAKmK6hVvtPC1WHvEI26xsorCSCsv2hu
tbItOcvduTJkv1dJ1GBYVgQz/0QNui97wW9IwQVc3zgk5ZpOA4/uT3WfZ8JyeaPAKVm01ztmbEDx
BjHDu6CufeCkCTwYwKa5pATaGXTIQsYTh4sPVfIFKcGqhOr+tRzDODCN/OA6YY9BVemOWfph7dhp
0K3UirwqgPOyPQGATmkCH213ArwLRiHAS5qlBL51gzOOG/OzpYCOR6b5wXpJVImlBQsmji/M5Jm2
ferf3iF61FndjsVJXFMZ6pDqRDDjkG1Aq2GOmFZsNT2OQnvgmd/OVw5DwBTjIKBauLTEHc59/bl1
qZKwtjuVDbIqzqjzgToLUwVtZanTaHu38C7VMg2Q5D6zUuly4AdvQeoJPjz52bvtDVRlgrtEjv81
ggDmO0VDtiVIwqY+776o0RCKh9WuVllj4Z4dAZ+gftlyF99D3QCIVbZXUEyaXmeW0gnlQIOdVaa4
Zg3iBbIK5KAY2HdWbcDqSsBPi+FEhigw5Uy0cH/Q2qOoGqIlipEuH5eAzVKzsh1GVvIzP2MHnjq2
K6eCcy/LDZrJnByW0g9Uj696t++AQ/8iyq49XbzHgM6fs+x/T5euGBwo8TWnAZoXFRJbz35LvuR2
z3SkN6SPdLQSTSn0sKx5R9cpycAqqBDlE9zmzXsHL5h56Kx1/YOCCYfoAa3y4R2YPwG4vO9sVcxz
dR8VI9KS5FQI82Q6VI9m9oNgtmP+xsCgiITALGorjHXGWdV+Jbr4DNes7zhLWZZxit6ITnb1Qcjc
NJeX412QvwmjLz9MzY2ahplLDVdZB848U/gmavOJfHNj+HqG/Nwh+rZZj3kZfH26PYn7ePlXozZH
FUfAW3GwALpJEOwoC68atPoGpANP77zip29sCG7d95GiK5hZ8HF4VWSPtwsbFHRN5T+pB0H77cvk
gWIzihhL6q22yAkT3sZLZkdbSLuGneq+qanIk5lcoyvH9cPe4qVx7uHW5JsZ5RCsLtGnpgUKrjcR
m1WmwYrSQrRZVR9C8KuSKlBuTNYZazEEN6EiSYsG7xwbAb65D3nH51UVZxW6f0aELx4L5eTE0Eau
nt79ICEmjg33emE19ofhNdJq0/e1HMHxsJXmaOtxE/h9EWNz3MP87HcB7IuKPUOeQdtJjZ8BHjWz
t3GsxQOwDiowIElv2Y7rp0EQ3PI7Y6/XxHuE3lS2zRMPKHLL8Ugf9jzQeIVMI7UDaIz2G87ZF+q/
HovXvy2kI47AL7aTCpEZr/3Urkr4PYlfsHeNLQVEwVleptNrYWdQxVEiB1UFWncJJXAkydeSJJGD
PtSJn4tnDUZAUtO2oJAEQKz15JRJXwhrxUL73NaZl1wOXhf7r5GyPbMps0zNTLmKJp3Vi7qLBiGR
1iTAiilNSaDNUJ/SZ7XmXDI/TxP7+cFExOusX4P5wNkjWMP3sJAhewYbW48ql9dYy8lDs6VKj7xa
gx6Ces1JAexazJ6ZqXBa+5472gj0YKjryfyThT4VIAA7hcZDrsA9kFDtVZUxvlAy6Ae6q0Ajw1zW
4T0dthLmBVoimmEyh90T35oZopH3fFCVoHdA5+UzSLhfesGcRpmWgOoHUo1mkntdvgLeYdpA+qna
41ND6cc2EfidrOsLP5DbjuwBqoto8ljmD3xmn3rvMmy47vpRdOkLJKD6g7fQqafZqB6BAljm8tDd
nfnu9htsz8x5h16JhbedP65pohX3BCRHa9tUrV1Ne0Ailv5g+D/DQXE8tOXUO7Av6WEo757BdhPV
hGGpYrfl1OTjGdvDIiuAG8mIRvBwa8fT9ESxzBmppzoteBLOxh+lZcj1uRqESXXdXkn04PdRKkPR
QTTf+aveNBneIpyRU4CgISUWsdrFv8hHeZsFSqEX1fxhrRWJJWTHWJg4h0vLpPg6ZRtC+ezKB0R2
xhYbUuClyp6tayP/lPT2dcd0+6P4bSi6mJC4f6YrC+q0YR7514vGArHrVuKWGjWUdV9YzYyIVjij
9shBlDaJ0D+69TGXpJUnYQoFHrfU9LPf93pJgqHEap8aL3B30dVMSSwU+UDp7/6gZitgrG35m4iy
3yksVWdoBxnxz4djk0oLJqvIhwAtz5HgqieHZYXattVZSYb5geiaWVleVUC9/HbxoIM6pmQ7WT0J
Waxa1ZxmqKB0YvXjuSoPgkzvOsSSnnay/eJ+Nf+ggFL4ZfsRtH7JlJmpiganPp9y6soT9lCZ0Jrq
SFn03DEz4QDmW7bHPzufm8J1Rf16liu5hyE1/m3gUWnRMwNHD9O2rwfXv4/iCkiZ8vX/8k5UHl6E
eyASWUZ7k8ElYb7a8B87CvuhJGOSnDZCObS/9iGGJ68/Uv2wT+tnSPSl5oUWE8ClN7E9tE2KiDOy
So+YpYFBYUNzFXzd1+OOlDXUxtFHKvYoJA7BE9AqMCTY+N14QazMCIPlAwCIM2ny/D3M/gYXDwL+
rICqzHS1+HYDwLb3z5hkcQ/J28zddUqBSWbQntnS1+AXYGjQYyNEESkVi4oQ22Hz+YQc1/tJVQyE
pa9uld/8OEj6wmv5wMnXmVwi3R84IsOzWJ9cswl90Cn0nz+60s6VknuJZ5VHKyqbgCz5/9ekDcet
s1zHS7CXUgZ0nODq+GqLmLj8ASRhhlDIhd46lTEP/opiT6r6T5mjskaUBiPmCn8iYrKOaZDduT2t
fhGDLsjpcfY4Nfof548Nrh/z9McG6r0GIPVST9B0lZ6DvEQ+N2fI9UnEVyMuRikXTn/hrCijBlTn
Tta2B2AJxf2r7mcg0wwlUYwXBLXbI0OpcaN9EH2gIpiUuXbSLKKW8cWxX3WuDbtDn84OKRaUGdAg
RNDeOfuU2WeSeNrwDd5GU15Zm3E5wGgXCbriTpRFahd/Ib4FTlrlpGJxU2w7I1BqnzWmIiB0BVVc
ea/QA67nTNnK4hziPtTIOvNYF+Tesvqi8sYp6zBs+Rn4A/QgkAsQIGjg4HiJsPRYYaGpdHNuuk/X
jVzhkoKE7qlmylCzpGnk+6w/rlEnViuGjGFm/KCDFgMWCrKWmOZttukqG8Xa4SSRLRVXbxJUZQo4
wdP1CmhBqI6h4CBgGEgX+50aXZQIOm54VPABKI6o7ZUDVgyzFbh+0Emn5wPX5Aq/HYh4I2rdtzMv
yaJYEb2kc3FDDBfXZejhQ0nPzDy563TY74js9U3GPUfr/Y/T/tT7aoMaXHk5ik6rtbEwW0T9zJKU
uLAtT5AtOCkytYDcTNRT82DP1/XBTTLbj611CB78jbYiUIOY6QFGcSQnQPY9zBV2hFvtXTWXcyMk
eoJu7Ky13s9Vrx4sFFBtgOHYfyja4WMqTc/ytLN15QQBSPd90cY7XnLwkYGVkU1eHxKOlVp1jaUg
+UY4HFKsGHwBbgOntkF0h0BUcHIhk6bis8mwqgs4gTFUPPd32OyLyfd8S6GjKujzXnXhDMSS9M58
zCKFv9B2G3n1P9ZkwAx8nEiS/lRBWHPnPRhUM0tM5r7jcclDumI9W6rjTk61WOu4eqONCQrGXiEJ
/BwUhwk6yUJe58Vs/0UgWXPYC59ycPsEeZFhrUYLsdUSIL2sZZu/bNII7WPJI7FsBhXE8uhezBg5
G8GFilNFb86hVy7//cdpUcsxkIr+lgOCcDxncy8oYhQxgqSMSaPPqG8dBjQdPwc4vY7CbG4AHTmc
kRcg+s+0qDQ6qXjciQO6XgGgczKLUDWywMP+aC5+PJGPNdJ2yK8qAhKqx2BFGWY3UoBjsqKv+pYY
QrAlcHg5X/CmY/jdpmC3i8chKSd6TD1GoGOZJdWoNExTDWOFWz61cYWv1zHgHwaVebicJw7NSkoM
TQQhfhvdvVGVQZriR6N6mBXkM4dLt8v+N0NR1RfAQwq46cNEeF/hpbsAZ9SgyYQrze8EzQhiteaB
VXuShP/VYWEEJLZ5qXkvwlImzaQUpt0UgAoO3jcLIpHccdZT3Jubg7xHSyDo6Ar3Y/sEA7Wo+4uo
qRGseKADakBJ6lq42Lu83EbMgEib4l2C3q5r5N+jOKhLmGf7p0pvwj0Wx9q5lOAUjIZ+RdenxrtI
3dAz30uFuRc9DSxz4keIrT0eW7lD0IN702WXKEmVOBSaot5m5XV0k2cB3Dt8wa9+KfJkQrVQz6v/
4XWRbECG3USdOsb0vbmZgc0K4G9LCLEtTxiuvmaUQm284CPplkWHBwRsDFVMOhW1VWscsy2dUagt
ymaTDBkxMTto6a+r7fINUIDSpKawcoB3XukAl4L+Q58s/72p48OvZEfYVPSK7BIID6/byKz66JoP
ykvfHbGm3qBgazwcF3AxkLI11wBrpCKFzjAioIME7LRBH3DvHnU70caLDea6H6PqAwPa1+ZLpm2B
jcsH02/f8ckbK1V+ItxggzHVxwl7m5ul//LIR9w1P9PQs2L0WhlFcm++zBIgINlHSkQ6KpbFAR86
0Djyi83V3DBOE99zV9+gKswC70FL1abB9qXgV+uCZWlubNgtpZjShqxQNiGrEJj5GNv4oVsYBZv9
j2nO4f/Q7Y3Zjd8276jpbZLfqNpJQmQT7XyodJgzLUc6CwvCRD8czgvRMeSpuEE8xo1ceoZwJbjQ
nCxFV5+cCGNMkZrvc/vJ/yhoORifbTLpjoPLHRueATUQ9YTNCPjzvxIDTBAh/R2+92L5Yb1h5EUc
BChrDK1Aid4fmSoKwwfwdNa3x/Tn47uEN6TLncw1h0+GF6bdTD/fFcu5zFj6iteoIubGUhMoLSDM
53p6JYE9m6nJ1cNtNQGujrH7YlPY0NB1zX688UpDC/eEh0w5eFRNFhz2LGW23/Y9mXrPrRNkoZ+W
vI4/OZuyCjTlHnxJ5UJ6nfhKK91iZ6fvh3xC01tKKrbTfv2XBa1ExYCQxyoy3Qhirpro4Jv0G3FA
EXROpAD5MjqoQLamMM3eovjU4LgJE0tlhMQhc9cT3IE4lws05kqYhN13D+CPFOmzDtQyVqKffl5h
aOTBY+gNWc9JrUtiv8PGmZ7li9tKK9EXhZM+MGZ49RBxXQerTBCwFDNf0jrTK6ERc0LcpKSgokWw
7CtktOVXES3oo+1OOo+yQmYhTzsz7Tplt4LVBCp+dhSzDfcz/rd3UzrjsA6H8e00HnvJHzKyM8vJ
jC6pEnngfFvLDIVbKf0sRtp3IY9w4N0u75cu+9UQPBwL/ezM/yg5jNqV9XZc09UJ6wEUQOn/1mb8
J+3D1gGwHL4mBfx71nVdqokZCwPvi+Vqd+0LrNNo5MP0h4+bHwlQC+E6s4CLkCTxqS29zh3NP1SU
1uWyZVADkUhysqXsTam82uv6fEEYPhmMCqBs/rFLcqmXUXcHPDNv1yJpFPaVxsDNGVvqacWOGaXI
1ecVLzUdJdNe7wBhJ83E9p7GYImeq4vQjLfPUGt894/lxG9S1d5mnsMwzvxkeVVE/WbbetVqbmyF
1Q/rMf0KQuF6qn+8c94iA9AuMX2yFNCVWWtdE3jerYCR4I4nF+RXpw/u4ltO3i4cTD2YkzQL8N06
cgIzj7rXXfLPbF4KEAE4ebe+Khz/beEK5fQctqWG9pcLMdzxik2/fnrP2yZ0maoJDgl/gAg9mVxl
aR5UCEfb1kqLls+BSXBHCDGzSwObcOvukA9C1vS+OwGSWzlL6/Q3AeGL4sSufs0yY2NnaF3OS9dA
95n8uQ9xCUvanZyBSUid8jlHyN5ABRVSojItfJcW/uPsA/5ZF3aRUlsloTsRx45BE4KvoSNcos0+
BUrm76fUuIPej4a+7u0P3Nm+jXuDoWkAprBgcyppMvh8fpIsrlsDNZGAtsr5DmjYIUMXlSwJU1TR
HjPgrPboJTHlFaYx1fQbVwZlIu5F5HakAD24qSrBAW/w+sGL3A3Z1/XuUm/xvuBYPNzQvvoaMO+s
WbvutD5rBEAzdTNOr+Fxeeh0peaOFLmIrBZcZG3K/Bl/biS2zrCnFXQyz9zXzq8N/6KXPYLcP44o
4Xd/ZT96XHMtD+1DvgWlPWA61ybT1yTgg7xLlIbJn+PUUV3MjhD7S34ru2AoG3aBpJl8w7I8+D8h
8HezEA0MF3YfXUO00l2sQRXazbVKxY1I7+y0EJIMgCj5O71QIqAAyZtmZGH/j4/YqRhiHeYw2wuL
gfoXieoXH3YDJB/mLPRFcnRAHRIbDjugZggrhQjdyBzmlZaunc2e8xlNzKhHSRsvqCst30CctaMA
1L+BLfgWYS7L+H5mbK6mYrwgJFXNfXFPI/DXRjfU7DhT9dTXFXS9ERk1ztODEtWsS+EGbcdyJF1q
EEjntK+8u784kIy2Ahuw6i/JkxeavhZKNIkbv8A/ovHvq0e5+aX431oMlN5amz5R6DPJDs/wOzJR
UB1pTwkIpPp7BxwaDb/k0Izf6sKPbgLKWMmtgjwc5Kbppp8Z+dH2I7qDYb1NDf4T2PUVzQY40X2c
KVlZ9UvBdPJz3I08HxSpzifcVZXClTkeHynKCvK63VDAMJ3BygbW3TC0CrFhbQTwiGLDPSFuck3B
lNOrxEH0USYWHgllapDFkfMSfmviDAilkHHMnhvm4+rIbZpCZ47WEImDlSFoW0Omirlq1cunvZoo
IOmeKM0QL8ekUs2i+FATfK2ZAWxoxRfdXbN2Mmk5N3aeAbZaDQ7eAmLV3+HRhyRKlKARvza87lI/
RbQ6BrNSSELsHZeiXXVCByuc6DkhZJ3BBmjxcsJoeeA/IOUnKmNS3Dwrun6tBWDD6wUo/5yvFaaV
F4s+6gj1BhxZZDRa1QxtfnKUPiVyZ2GLeS5YgRalZDBe8Fij4xFxwBwXvkxn/0AMCXdWgE0gxHIQ
ZFIlGdnEoNiUBefZoWS9B6K99Cp6v+HGknjiZwX2M2XpQGJArW1flXtFcD4qZUGycpJat9B/Y7Or
hGS+Gow4At22RE+VVfw1Q0q1WyJbheECQtuwu5dr02SKGnql033B21r+XE6phdGSroGhLN4UsLVL
nZnXBlySE57UPoTAT7voJoveNDUtt/TGPdWvIHcerbYfyE4h04x4M8On7uIwxt+lUuhLOEkRlTtg
mEB2vVaDthnevocyjRd5nmjJtLYCUxaC2hKAdoYUDtXS+6KZkPbtUWmwpF5R8O7B4hoK0p87Rv+l
kDNdVUSXVl31tiEroP+kC7oEUvJAaAUi5PHRJzi357cJ2e7nisV86FGwp31L1CzGh363F9nJ2HyG
SMHVn/GwCZtBAaGZZwi8pW8oW7OqtinNzSMh7V+5Yj5vngBHyYUsPBSe6KdkQMkWOR0x1Z5Wvl+D
OsoIUDTAdmCv2+TbQqHQylozGDaKmR6zQSpkVr2iUU3oS3EcKps1x4ZgWSL8LcA2jwAByzW3OmrB
vF/2IIb8n82U6AXbtDfSQz/x5FcdZmQ4QjdAjQYIz2BoS4Zs3b2R1+KkOSARnGPXax24oOxF3Inj
dEyj8SCLHbhO+jQ2YYZYoEYl+qLUQW+v/f5xkl9kBSHZ1w0L/7HW3sjH2W4HPLZ9QLdZqV3eZvEn
jsHB9Lxvu/xKSwF7RDkWf7ESZriZ0C8eNDENMuetr8NiOuhmZbXrrtGgANeA4y1jBJ+T7+Sys1Vf
PYxvNcXUTwCj1v3Bezqk/gx990cfUaMZsE0PQULTnVDj1TNrqyMPHludhlE0kGiLCrR7ufDphSyC
kCSyLoBpWmLsvp7vqb9QwT6VpcPHX5PtrAvQRMD6Z9zx4jhnnOq4cZSfczMHkxwTem6i7nss4TBY
zxZHUP3oL2nCW4urMKFObJCKQeEUQtVmcEgEkSj2sM9UC8tTyC6vRI31YdtgshchQp0QrIoh5OiN
cmR3iLgoOhYqXdvPassxCYxmxP1PYgHjjZjrl86ct3nc8+8NDIEA6IZqYDmF6/xth0/H1NKTGGgY
1E2c9/0iaOKYpXu5BgOBY36BWu+t9X8frL/sH0WDIbgn1aoCMdo6tJTV8IS18TZX0bY4vNXh26GM
8EGPgEIX0vj29qCcSposp9vwC8mE5njBnUNEodKdP5k2rhlK9P0RvjjT8CYzDTxHvit4LirtAFrS
Ct1/B2w26jvSKD7E1IyBGSraVFdb/Ozd7ePsBky7yQdEioD/CnAD+r5ANd4jw5NnKCEh2WqKtYRu
XY+VNZpy3tuMxBguN/6ATHpKK+yAw/ykrTWdEapt8rWLXxJUgYMbj9oZpSKXzNgh1VeNs6N8NViQ
3f3MhNbhO/3bbomywKcaScYGo2JSi34LcvL0h+ZG/VFSNcph+816JI8uMNCPR3VrlxX4WoXpLQKf
+6K+GZ601QzDOll4BL67k0pl5SYPVRvrMaH2l2rjCnY8mVmR5OgTRT5OXLl/wZS/j2JUxWr3UYWQ
l41Fw3LXSorsfRx1UVbcsbH5dv0671nVtfSP6P5JYf4/jamZnPr3sHGOC3X29W0tpxNKn4HXqvW9
brOPe6OCZGTi4/fEvKnM2QKUHZeNjeimfj72Jw889Aea4k8Kg3VAMzp4Yvw0VNYHqHR3zoeW8FCi
lXK+xrtOpzWGTDkRU6+aCJw5JRsiWhh+RAWliatH8zBJ88NafBGsxNtY0Ck2/3dYcAf1PJwAbywZ
Yh35O7ZY5kN+PKUt+v/xk5+49bNEBxmMtaBf9dJ5/hd3/rmC+E5111jeYWplC9Vu8Uo4ppzGpkx8
CjH9Pma1MDDyvCluLnuiH7JA1PucsB0XYsbAbmo2fwAjUBIqOC2rzPcPkMmSTU53E+2aUqIdUxUf
0fUoMbCtIitzRs2SY8gZ36j01gqazMJvHwbsuKlFmjSTxRzdV45Y/n6YTjq/t+bDdzhHo0vqWWv1
mw5N7RiroBpIxBVwaOQfGlyhz5XfMy/PTm17E6ImFWqU4cecPx7Y/13TBWAAgqsPhBdDUCjq70x4
5AdydsubvIDq3KoTZywY3f/GuPhs/mwBtPjPnBeo/f7XjzvNR+jsW/yimthNf3qoMnYJZUzyROHQ
cV4F1PPO6bApgFQZKMnR0waP+/1R5I+cwQdiNGmhnU+AD+BA42aWnBtGhk9En63zpYG+Ptb6+/T2
o82bCFyqvg3pcnnP52QlZ5go3VNwNAMMb+dBSsrK3W6XgZ+F38bzhDWpgoKo/u5AtpLvIlvprEAx
h6sTJwNcG/qBTeJco1rcID96M6Q2/VN84R1n4boa8qx4GX/A0TYLrKKRA5WD3J6/0Yrqnp38KL/z
dcREwAlY8jc2t4XLSTx2waQu6Sj9TWo8ll8idgHukUw4Wrmzal7wdXjKJcHMpLo/EgxmhbvSw4AB
cxxZRP4vlkE7982wF7wwUdHKPLXlD5GGenvKynvUMQ/ZgpEwpezjOeXi9lXMuBH8VvsXoAML29v7
OMuLnCOO5EorQzs8U6Y6CGBm5ixJt60l9nYG6BdLcUjRMSAxzF4pJbpa5BF5VXtW1z1pCSTseAcI
Q6pGXsnXp4brI6rDgVHj1a0wAgOYy+SoyA6xpaQJ+rSGcmXoo6HQkc+aFTfOn+jNm/ZaVFd3INzD
UnR9UjyyaqkKJ4IYL/u80bWq8ofqKu8K9GzAeb9s9d+tgcp1eMIJJSbOJGV3N1Ta29nkgyRkPr+9
45U/yUxm2rrH3I3XPwb+slmKBZ8QxXU2Mfurnaj0cDYMgsaJDe1eoavMrrf0s61RIf1l7EYpwrcQ
SWyUNqP4uvMWCziaJX9mbagNoy6rqa/I4om/QQ+u6x1UfWk8znE6P+hejpHZSW/3YxZn6VptlStz
9FHo0S8QIXjP6A9Q7CNV/2l+etaxLOT4J2hmUbD42AURzzjn5wnmNiugEf/YxZuPEFEoWAJlFMTE
rexa8JJAZO1p2V+z+STIKT1aI++KUeBKD01E3lKAzGVXB8toxLIBtAejNg21r9/365J1JPqrfjKK
RjWQWB6B6AdNeVYmmcQWnzckj/mmqUScF3TC7o+qMvKPMKgOIfvBm/0muZcUSVyNPpm9GJl4r3vQ
NhBthd36Rsp16exQDwPfzjla0g2M0iz6K5JjTS/eW3BCLrg2DJPc70OvRlXE1U8F2qCJ+Iqel7JW
gG9alhQ9bfZKgqsV586PdKsOLxYsBArw1do9INHR1gc/zl6vueHG8Co605167D+q80028mrNUTcZ
QNnedRc5L4anW85tL/X7hmUwiz69SSKyX2diEMNoYCKkzShMOTVNwUmanofGT4pSKjwfVWXWsXMq
7DCs5uHmRLkdWoNnH65LNzJsOVZ4Jn4hdyj3lAd5RT6l952d75B3Hhm99dJEixrFaOv+40F0p16/
dWsjJH9XIXlOYQndVMSkUwG4xERWQEXUQeHrLd0lWmyWjUblZkGMnI0kkow9wK4OL33oKojQI7GG
e+s+PRohnDtngqtxgM30+2SAjTtb1D3o8nQvW6K8GD6zdCG9c+hSP+KKqnIM6DfvrsytuJfIY+FA
WgYWlRGt4J94vScMIyqcz0KvWdM+EW26xDeQHU/Vz+8vydxgDfz/lciEjkNqVE1byXnbhdPPS4Uc
Ju0amSar+d/hlyaq5YqKv7C2Sr/1oeni9w7OKVeb61JhqVVg3w4OR1Nev7TNUMLVUbAbx0Dua4I6
aciM86uT/OCV6Q9b47Y+6xR9TqWtgfogBsfzfeDQNI+gANHzOw52jKPjnn2nNHyHhtbSAhn0sU+9
kM5rVHZcoVl2TgAySArhGF2UfhYvpsjYfhbWIVAvy2O9LK3R2cu/4blX4oaS6G8CPfvtrXc4Wk4y
YWfTvlxv1cG79DeZSU9+BhU1pbiNJPbF1+WIe4Tca0/spLj1KPiylOEou4yQZbL8NTDyJsu0lU2b
wWmbQgwqCC4jEIfWsvX6jAXd76L60q+hWmIUeo0mdWrIgGa73l5bQX/z/9xg8t+L9jm1qAMaeOmi
tFLZspbp5bciFVv754rIPd/NxX55ad9AzFXNyhUoQd1T6idbFZacyD5Fg7I+mLecRCfH6lT1em7N
sHy0JgSdlQwrdcNJg+CT6xVYcDuIrIu3gX7/XqIlO+hgj1vL8QFyfSqn0h7F1kbFAySjRtDXE0Mt
bPwk/NFqAEB55Q4/Q4f9aHeiA38IL7cFOTHdZm39sjFQT1CUg+bZi+6BU6XIipV/gmL9kBc6ffwI
2ApXesZnQUgiujEbRlnErGbzK93TaiTEQ6EwRAuV+UPoVmRj/Am5J8EkY74cFgx8MRm3cNfTGHiW
mRdjwjP0vNWV89P9hK8UFsWgREEzTv1dyNI0EoB0HJ07ujLaCDUv8IiF9vWPgG3orgfbBPI74rGS
2Mwhh3fdJDdwPSSP4OjbSIwuF6mr2NKUzrQ6KX2ryy1QMjBb/Cnf6mir2BeOGSZ03yy2oh8WMV4B
HtEb7E+KguLoqymmVBJF9YpmmHdynsrlydv2gezp84avygaV/jYJquG/4e5wHzZh8rg3Jb4mtjcE
M10B9ePP1OaSyxXRQ2bAZ9vLUIAeceLnxGBK1lCdWk/9JXEkJpFkSwFsgNd3iaValDS03e+GD8hp
Haro6Ts1Fs1OCrPzi0VURLWStqMU1RQ3zYWyKwkkXmy8W1Lx78bV5ROBswUqUqmZzvDURAYevHgQ
z6kSgkKStokMuhrkfNqbj3jmDNkZeSfiWbiyGJGyxZWN99sNlTaqgCXhdugKIgdb0ftxnwipQv65
5s/M2Arqfe8X1uKBS8dJRXDWlqMBZP/KigK2Q1rJ+cI8EFJ+sEh3hYIzkb+atqO1v/HkJHefA767
r+FEIPzO31FBh1quCou8kLTAVMrPaw1DtgxSKLGhHxpE6hw8c0Sr4lh/WHgSK37ylgeAnO61iABn
Q1SbVxdjClB83juqVId41dpYG02WPU5HWsj2nkjdVuOrAG723h5nr0q593TbF9WTtxQElXXD+kfa
r2vPX07ym3R9cfBcBR7BWkDWunyJXH+WOLTo2VgeDgcXWC0ldT2IJpO4nTcHG4ilgS4kiSB5GjEi
afRwn2EeqXU1F0MXoPqXk4jvvcX40WtAYxXZx+58v8rVJD5u0I5UqpthHNrI4kIb5NGv6xuXesWa
awDuG7sWzXBnH8B1Sdj48nxatH620rJr9TS6/4WnvE0u5+vJyxMshcNw9w9wDVG5LKVjZcNM9cXg
eRYqVsLNN3dW6BFeOwHW7AO30+pHtHY5UsDbKcDhM3jEw6dMJhfPZfxqPotWKgzMO2GWOruMLsAo
kJ5ciUVJUVyCywOD/vAlUqHOIKpvwmeeTc4pE4i/GtQrGSgPZN07pWzajj0rsdvZ5viMs6nl/ZAh
zxpbDWqtqER/V/Vz22/i0Q4LX6Htpeu+PpFY34W22nU8Lo8kqplxeT5AtfUOQshSVuk5YiI/YJ0X
vmzjbIPE1roZ4JxUfll0KHTKo3i+B6x2VencfkUFN5lrjyT2WkTu+iKL6Jl5oq2espJfQuV+1cNQ
MsUxTlfKdUbVmZDwhO5CNrUli6RVk6xPyr/GW7peaoZmWGMETfRDchdHMQlc5Xq7XPwLcmD5MV4n
hpS1HFicafE9OuPgNwNF/dPjQrk2rULABQCL8e5zBv4PLupimOcPjYYolPxKR20yxxgkMBnxPuAX
2j7KycXUSpZBP/EqUNsehGwnjTloIJqO0JXYGyP9GQVNP02t1oS6KwBrJDNU6xc6u47GsG+T/3sJ
TBYfWYFvTfYdpst+ptPYV/eSe3y/LXMZsCD04XtGQTY4Hb3x/1LxdAuJeTTh2On6B1ecNt9b9Bc7
GLiXv7nU0XYQmkRGu1tzplMrv8EZ0eTG4tBRPXB5n1scAVmyP18VkIaBxnCYwoT3NcVctm5t6KbL
PspqRsiBUWvC566tRAyU96Zr4C66Bjxan2b7fjsXfm2GCfrXl1h9KHqEEXKibff5MRb398gWVcOY
HD76uqkka9Zx+llvmLSx5VBk1AKKxwET8v2IRTKIr5Ytcg/MBSNjlfYz4MI2U5180Xe7HpgB5V2a
VIg+g7Z3/4ROFoSiVrdhszn3rjjT5N9qAer9DNDG8lIJ1TqjA25dzDDD7PsaaDLGbzDWQlvyMcI6
JkgZjXJSKq2gBKmuISWjLfgz9spXJFrHpa6FSGaKYPHEZZ2w71eH7DyGZ5gYZAuYbupeFV+8QtNw
BClfA6xsWBukDY6E6I3ej1O70RelkFM36Ea1MzOBG8AKzH21EYNVkdjIZKLOTqujtb/2no50qHa9
bvtajEzTui0gVz9/pxXtTn5FRQ9fe+Ugl5h3sXqakmQcGH6er15ZA2UcSXgMV7xDH/p1dwD8X+Pr
rTIQgigB4A8SyUb4jQ4MYeRdn5N74Y1r7aTEgyBht7vn52JCB0dDR4/zTRJrRSuENuUbh95MBbpj
uxTmJp0J39UjdIGmrr/jANuGxOITyO3YVPMxWRlSF1oqdg/i6DElMd37CihRoRl1PfME4LwEjWSu
Kbv5fOAE3Z3hE1hHs9VfleSdbbk4InWt1Qaz1vHqZVhIqQYB7xH05ovALu6z4tWXnyEOTYBoWtTv
iYtSF2aXzunSd7qKEtmEQAhKlS9MmQLlancSU3/PBl1XEbBcPqBpGXXMbeqnc6FopbSCJMFUAj1j
EIOZji9vIZhTC98cu8SMfCeEwVCnbBWfZZe4pYMg2VP6yUpHQl7+6agu1SIWMneqRQcIL/GUzqMJ
lmup8VUo5MpMwAzC0eY2LZecwQRJNh8cRsjl3SqfAATqDuKoJyMZrj2fAtlwlwka8IhNRWmf7YK5
I8sgIrXo1X+S5IK+4nSg7It2DfJOLKCdNjQhiuYDO2ZV8Yu3+I6ZkPJV4uhtVvNG+p1/HZMXfUus
F7kTxuHUmwIV3pZzQwq24HOxlD58BdBqMS6/+ux2sBu78HfMPg7hD6xPIAcRomr6ZDaTtVBRT9r6
a5ePjCW2v1pJkctYKNKxo/op67zi2aVZTXYMTCix+6iW/I2Y5gmMrLJAk1czyE1O2QMUzx8mvQS8
mvv43A5XiyOIzzE7sBJOXrVtEY6zXmVtdrSilo4oZcwy2Pg2rlSru0IiTgckuESNGghOuXJRHLDZ
sSktTmFAWYiLBUuiuulxi4m9Q4E1ysRAS3HPaOsehTRkxHeVe0AlzTkjykBbj1eTq3LCWATJMJ9i
ZAA1FAWjiA2AjubZRlRPA3pUofqPHIsel4csSts5FEBg02hQtfEbsmML5YCy6jrVzpM8fMXIdBna
/ayFktrwWGxiEOvrFpI4/bx7OimxIO7e0m7O0xX5cMzGLXNrd/hXg9kbjy4Jr8oP0TN5yjIrBOY7
LfdqWvVs4ph230QafDTJYSC6tVcq8reP5aC1uov5vpfltTMDq5ZOkK5z8F/gI/Il6jc5DtUU3pmt
SxV+vsJ/6r1hlz5BmC8qSCIlPzj875iSPsXFZ64DUn9s23FfpYDRYzRlIbpUI/k5qwPWqNZDu1RU
dKWzqDU/n+c9GtcDhaIuQPzDkgyOw3EQsnNUiAO8BPaoLNntfN8hchXwuCLBGBBkpekINPa0ytSl
bk6kLJT5cE8gcwUPpFoaoPb/Gj8uIMI5YC2Hh8Us/x8qaA2IRDTQqrfTvWQ2NyfC/njmUeaisy/7
IdOWmUvrmf2fCIpnwslCYwXRMq7y4A8wPSWzXVzpzYaUzSWi763bDicXR17zTGuEhdNOtwv24f9S
8SRbAPUVoszEYp8oa6OiFBba7KLwcl749O7ADj31DB3yzIdfU+qR8b1v+7VZ/Oy/Xtwd+Qb2SAy8
TGTfr2UhgmADNFHy2kOTYT6yLJyt4ceRW/pK/pUxFxQzv36qTCHwhMlIo72rRMdv1v01JECuz8iL
07RB1KlX1q053xNLw3or6kl+WWCMy1upuyNqhar5wdcKqldytnRqYt3VFZrwBZXw8dfOWTt0FOJ1
/DIFtv5Bs2FEhnZok2304V8ThRGZvRJTOBckwsE35ZNbeRvrxnRwcz1HvmY3nlReVxB+HVQtdbQ6
J8adHSfufIJKcVdEGE6ejB8EuOb9bswqlnPghgijtCODuwa7LY1MHWa6ZccYg783a1wYa9vP09Qn
fKHCNn6fUqnFknDMEM9AJTIeAgVg3MFnWxqnodqynbpR9O9hphzlpsS77ThXq3guGLLGcZfQpopZ
0Kxe6lVljFx1Lefc9tZ5gDnCyKCkdjS7LEOtrLaF+rOPxJgIjKZ202EPQ9WRU3xioInC7yEa/tsj
P0/h428ZSFWGoC+y43erl7hHRPyGBdT6q1F40mufifGtWeEHTVKldFpwo53/v/WhFtOltChux3tu
eOuTSjaoTb9clbtBa97ImQP0NLffpI/USpXabq5vHZt4w6EKuyP0jPQOt4JIJiWlL0610AHLLgkX
MH8Tfl+NzqhbGQbzhIFMLhgOjyiKWWEPDASAgYXHxPXxht97z9UNLYZRJuvTvryajMSt0dPneCbh
1sKbjR1vErI8XzZi8SVxvDDkPwCNk67a90z9MAgopMfqPxg99f7geOKlHXtZHCo9Mx5Ue22wkqJx
ICQuprxjycYr7oy3WuKTOZxSLK4UNPS7yqcBBPTCUGYC2U1FMA+DsVSwcOuSWtkeU+XngqnWzfQA
8wCz33CrNTQAv9vXMhJPCIlFI5FSW8ZZY1/qpSYRze6ezzBhtcfZfRt1UEiIuM8ikKfmRCb/TSqz
jv6ne4eEKAI7tQAm/JmKLiYrZXPNx6P3VUoTAoU5/VeKP17xiu7RJcbTu9NEKgmjtLOgGIH90bE9
9Itsqk2q0ZkQ65Oa/+Oea/SDmKTHKjIq4HFVrmixmVtIrcc8/67fG2fY3qBkFR2xhvFhShj6ALu8
Vgu+i73Dz+9jacyoUDQ/3+Z42HrlnRbqBX73mOgXVv2pcp35tq6V/sbW+mFD5rhv44r/Ltqn3MxC
XpVJVyBoo6jV+KtfVPJxz04oZdetZpA1/ujBzH0LC5IcgCbXkgm/anof4ScYaADKj9S1T/2HPK4y
YKwasKnyEC9SUsEwGd0WINO6wYe5tC24inoiOMpxFOqgnzIBxQfQ53f/6HA82A+ngRVHIMWIXItH
aluKNmqVMuCSIldECYNE0TRjFU6gwAkAUxu6EiMfhjeFQ8DmlAZlNA1p1BzjpjN+eyzXeaIxPnqJ
6NuHW18KrgqVhfZNt3u6hOpEe0UYnsMLbFlk3vTHwrM6ONBJ2SLg2wEI8LUKqQWXu5JGFRMDTmrY
663+cwq//ILQBMbfCT8ecQk8L36nr6HvY2c3qE+ypxoea3Mg6knsF/PCHkxW7OjWszsJ62UN4p7t
AzXsGj7vD6BMG/zHJt+F33NFDvskGjgDyxwGB9FtOusniTP5ZnjdZh/uR26u7Mamfjg/xqR0PrXw
SIzNso6RoXS5M7r0DHnN5Aq0vCiepd/v6Zs38t0YEadpPGDT3d1hZTlnX5R+jD1F1BbBWbt3BOua
C4UEHYHf6Y7oX+wSbY28WoTFNPcuorxPhoezV8nHAbqSJJKl/zin5a5gdk5b9f7o+qEsYbfJua+l
gDRfmcWil16akXzo1S3vu6JryVAR20+osL99calwso1QdCbVRhKlShCACVJZvCZ0JHQAZqlOnWvp
WVxmfL+J1QRh2nvK1EzkrRHnlPd9lEMl+Jp1/rtBUP+Zq2EQgCucseakrqIKe2BjUDqksW5mmt6G
FU0vw8U8189rEtWFaDKlts/gOE3JWra2//Et6sZzGJPg6UHuwoBD3y1gRoJCTZN2QJVvE4OjDZu/
khQEiLLaQk+Yuk75r8K6rve7I++XGq0aekUUrTH+rz06Jb+es4F4gaiUfDEL+x+tHT8UY9EfJb13
8sZyN2U3GhONnDkEGvWWtF6nSoAXIoL1wBw3owdtdc+0+l/mXuc0UAWFbGWB/edsdxBppxMJTFSr
CbkLToLr4dhmvEhf+3DLEk17W+ZhUrauOxBFdf27h/NFNtE5+vXCzav/WYenIK3ESCNJTpUVEekr
fr2zluLhthJp4lpk/FzoG+voM9IwXA2Mi+krGsQtavoU5ZQH1kCMnPQhd4ji8g/ZFT9Yb4aVuk87
kAa2sTiPbWlBpPBn3D4kM2tflPZPIyAzXYbNK1faenBxG5p3neiTI8qBWDS/tRoNieMP3s96NTjT
G/9q3usx9jHBeYBNjsHh8aYrpCuP+lDkqlvNIYxaOxItqKqj8cc4I6FjQPFBWw2OUmJIcw54Ticc
jAkph0ACbUOAW3YC75dOGrQJCXWSrSks2XT/oZYGzm0WwIbTLQ1JGiHJzg29EbXgLE4m8U/E78Cn
8AJCOX4bue5OOe4TKiD2IezEeJDrOoycw9+ubDV+4VlXo8sxw4JDlXccs/s7d4IyjM8/0DGFtjpQ
RZPPRtlQoFnrGJy8wStIxtyliNTVAlesokmmRuEdm8UIXSeeA5AX5Epp4N9Ac1S0qT86MkJYV6hC
FAS/ZkK6FTBucSwvY5zeS2sHKcX09vLuDz2GKH+TXU6mE7uHQUz1+5pnfd0yYHXdARrMD6JCRnuS
O0SbhElAVGa/q9PqPKF69i3zhPmHJ3R9AWgYUPdhLxfctatRDqKbB9gjcUGAH3/+5NfeJMDw1aNm
e7gfF3+IB5gw9go93dJx/WFKCPcuPFaR0KLPkxt5s/htExSsz/MXoHe/JtpsQRU5+B+4ZOcu58Lf
QkMoZjc1E7is28ecUMrWsyn+PRuYwvxt5dvyOhexvWh8fUstIof5noyYsWAgCKnPOvYxUF9YyC+8
za0JCcD6U0voNGdOM+L8bYxkjbqlzN/3he0TrchmHOksPWvP7XHU6+w0Ax8veTF8m5+WLcOYjibA
khubPYS+T1DsZ/NCr2BPKLQFGOGqKkdeo3H1CORCDliinwlrSQuS/wPgzl/yUuN+7BusJiQuI9Ma
0YqtjabXFCf7tZ7EEW+0q9gq5BSNVK/nROi+f2stTXEc7IpmlMal9QtGmk+YfsCubdEeaRTuTGob
Dm+8CTseVsS5ixH73Oz98K5Mj9WKFWvMY/24DRKCnVqb7hv/1/YzAOGZ6gPB8AdkFZNxYuTpyl3U
1CC7+t4kjlK2zccgG2NThODw9pJlWUmkxhjsQXCPYnp10iZSl1KIuUkzKWdrGrqAiSHPh1NjuRMW
11yLeRuN8ECImFhsnbz/k3iR/N4zzct22qce1n80cRG+f1Ho535skC5OKPlBVCrEkfU4m5vhnIsQ
X1aYmzqS+O+y+uAZHt5hv8D4WpJKgmyazbwmyQE5XkWlUpophFPEbM/cQu7qyUWrAhRXzJ2FLjjm
T5U8uEyxE4CA00JOkv5+WxC2n5HcTMzGEOkVssPQxogAcSbdRe6B0m6JfEBnfr5CgTYqpXlab7Cw
8JheRBs1HTtJXEYIZHvdT4cS3fR/JvVkxo9PGnyHKHfdYHtyLOoniepA0g33WsMoB6c12Fkjin+S
VuL+XvaStwbGEs80Dza0OF8ozKEQdPhzaklUEhgM0IzDUDT3rf8sbCp+028+H8y0jg/XGKaksQYi
t112Re4FevX4QKTXLqWlsPCWyGVh0JePBM2UXgQXHug39Ott+iKFG7bFZbqBIkI96Hgs+aXDjVCL
CqHuy30E+te/HlPNM6MRGIOW2erQ8W3mTClZBw34td/m0zGVzdRTE8qgEeWa4Sd8eJq7dwQ0QVQq
EVLJbx8zLdxUttqLa6UtGkDdI/M2aY8d29M3IUlwei8xsp7Fesf4+7otLlRmcUknf54Pw+Zr4y4Y
oh8HDhgRBH3Xr6GgOHN1ZPAkyavksrd5nI524qK08QPopSp2qfNbUaoSGojUE55kdA56oIaBMj6n
5+joOJ9eSIg1NNxlKyCd0DCN62f0ap6+sdWUsoEA+yV7xStOZaa7d9d7pAb844kLAaY80I2/45cK
v+XmOYVU3QpvHJqctXwJVPEElEvVc2qUJTjRIPqHE/+eYVzSHLzooTQKPcYhjmJD9kZN0i811GQV
+7ovcOtcRzPCfU4SmOsiupfoYb8lvuZ18JV5em4j5Ed6Gy6aZ0WgeNyg66TRRlLtDVRGlTmRvbi/
2febuW4byXfp00Xk2d/yAEtYHD7TwljtzYUfUYf+q6zIVmTNxigHCBUgmWlk6Q2CawUCSdNZrlqX
+lM9MQVbkMc3gkPoF/+QPpLaJBb2Cu2XmHIkt4P+Ne7OEmihlpC4iXwy9kbHqdHaDZpRfiV2Oht5
6Dlw3j3xPCSueHMLW0hoXjt36eKQ8G3DjwXDRvsWPW6x7B+Ob4bGIHCNuUNP+KQ5Ojorx+6ZH/WM
9PWaQsGdrvQ/24uz3m5l5Wahf4qhSBFKdr0+YQ7FcpGNvxFhi7QIDf7cHxQUyMAwggfJg4aC3/F3
2JUrdTM8i6d1GIKa/g3vXF46/47h5QuYa4PmEVk9xVpXbUxB54bmj4PfZebzyLCVzrTTbY3r0nnv
o+ORIOJz9A52hUsuU9qgNkh/c0qlT1TsxyDNt2FM+75ojoodgfnRhHGl3/7XpT9P+EoGh76+bzRU
tzuqJ9GyqLcXOiI8Q4WnsHyZvVieOp50gltnyi9L9G+1TUJzAsC86iLUo8shIZuHSpXIjk4zijNt
R11h5BIvLBgAPa325tHdvg3uVYcM7fK3d859nwxe+KasjIeb4ZQRZQ1ky8HZOIsqhFrx2YA5olFY
wdB8KeCYJHoMytzSbQj0umR7bTriN1dmUCZCUOiBs3vxiOD3mDw5EDkRarqfHuHc5r4oxngYi98z
Axu3+ksT3UUMoepNEFaM9NgWtobZLqr89WpGZgppkXa+Ib1VFxg5f1PEqMY5QNaeaHY4oP5t+i2n
T+NkHKuVoc2Z8NZIymuKq9DxT9uMw6UvJatyco65xOJ7KeMUSE4x5B/MPfSiSJg/k1JUYHXHARCj
9+hP2QACxn2iR2DEiw9PVAweEYsNvZ89FhSrUbifIwjeqRmMCitY8187UHsqix9hpzBXQ5+R2DOc
NYuHF94RngSHZblMneHb6dlGXPLaaiOTQfiC8eNR56TvMBh3sYE7KkY9oilzEcy6oQ5takWtDicn
bReO+nv7c9h4Oxji4jsOygq8kwxwr93YEmkb0IVmdNMjtBBTGTFBFIg2BLOYvo2CT0w4XzCalaiW
/IQY3gs5mL+vODlKWkqFF+c6pCP0zvdiYxnA0rUSnS1R1l9ZgR8DxC9bTcslV5oXOWIMCze3xO/g
fgwAGT6K2ZmJP0ZWwj/rlRXrSOPfuK8oW6ORDymy7kMYtb1BQlpuKKxPKg/3il2G03KHsZ+yb6jR
hxShUPkzcMu3b38w8ad3iRAw+s+KS5pep6NtnYanp3AqSx4cl2l7U5VZVyJpopwin404pL+M77vq
0zE9zR7Bd7QHEOoUswLKWeXaL90nqnF2hKlmcSk+hsP10FD6n0oVxL4wzopAK/fYkzNOY9jz5yVz
LdkQS931Nz8I159S/736gSIuZYdDJGldCXqiKRGk6woOdeBXcgF8MhE8mVyWOtqdhk7yAHRarE9t
QRuSI/xsSK0sDHjG4xLeAA1nAH+7HSH9cBw44wzGXvgrTaYGN/MPT8+iHIFRbKXcHXtof/6ieEpT
bBDX+cHgJR0aFFKD3dE5kUx3O4gbcpNKCZGTBkor4Xt60G6omjXjL8zAAP1EoKye6XSw0NbxaE1X
gWD74WqbGZHp+XkjIrQ5JpLlX3NfxCoWGxk/675ktq4MbD4XmTzzcdqkqCq4rvjqoHud62by6JHn
+Gt05KsZhzWOlrWY/B4k8vFb+0WOSlXXwOKSBOZEXAiOD4gbe15CdEkoQZhyZB19R7eDYZnDUxSI
mrk25Fmxg+Iw3nZIixfgRceKnc7TwqiSMfd1N1M6J+dHCcEc8AgvbHbj261AOEPhkWXxXPvlk+Jd
8FaU4AlJ0uvJBmB00Ermj8XgyoS/0oY939FcvFBMEzlVphBZYEaZD0CXzVimPMTikeOFl09hgDdh
m89hY/ysgXaKKo0c3eoKIzwSagjjMSpm1j0m1Uis1pey2EKxePTCV30926EW8e2NvBe863jpJRYN
UHhHKAfHRuvwcft55jScQEnyAq8fO0OYF5U+B4tNxUFNZF6fLJt1GLbCD9kDbeFzZnLTetE4OS+0
gOxggjf2XarjQ4xJ7MyH8BU+3KpjaJXUleeuTsaD5bqsAeypCMjPVBXk3k0cz4mKO7Pz4t0POSai
VPMzlUpcLhOLl5l6UdAoe8eA3YVzKfaDD8Cz24KAEJyHaR5YgCvCHMDpIS3Ara6oorLRkxTeGL0t
9D8Yup82jIbwzHGdBOLuQ35jGBcC5+PcNwLMH0HXLTXmS6xvNGuVcbSFnVzsQiy2ZEfc1Vz9gDyJ
yihE35iAh6icJahmAkgktemM85SAILxZPffTjbxnSkLoG9kuoGzpLv24jT6WRqOAWRy8DgZRzxn6
fYMO8cGJguuuR5PwhEt1fz3W1IB+Dqhg4PHl2+14sJcJqNl2sfY2UevPY07RI2XdFvS7RfPKB7NE
CoI5oH/uMepQHdG2bc7Z9jGOaNMl4jhp0Q47KVGU5SuDu09G0IgnnMsJVWimw6G9XaEB3pHyGF2f
y7ixE2Iqv4PLddGzAX00QmEMPg8T/i0mXv/F2F3DQ0EdcLqXclaeCsTqAFurKetKPHQanuKXdSY/
0fTLtRnB7sHurynAoR08AnJ0YUq7dBKQsQNqWV5vGSm03glG2mE7NOxupJjlZZWJswDXhTBm/qdW
0AnIbgkd4+/I/qQIMa6nlqHCDvZ3gl6nnX7qOnNnIKlmJ9JjziT/IHM4RcYgBJJZt0fU0My1gT5m
myxCgi67tyq5v6l5YPg/OVcFjat4hE1si70Hazrv4S6ETU05Th//5mc5/3+Ik5WbhBqaaE1+ipwh
VEmoeYgSjcO/bDv0ZAvzNXeM/zRCOfvY0OjFOG5DLdzQHEFpZAWdcL/tFkDTZDQPmQH1RjXRwmU+
QuZio2x/YfxsbCoB/ppuDxu/b71DZSku1prNhlqnZq5QhPlM2vT+MzOI0PtV6aCSC0ipExWVGNn5
UCTerYKi3pQmvYXdllPdSX509tX/sOruqGsvZxX1nFkxJdzYfRpRuEiZJUhQ9Bes5ixk2s8DWg4K
XUbTm84IPp0qO4B+yXccSCDgS+QhVrkqPWbdugJEG8kA8QsX+uBvBpI0cMt53wCIlEsY/dKbQV+7
jE8TnzpR1RmSPyT/m64Vo0fMNrXo44866XmKfYx17P3atyYjjxymg/W6UhKfmSR62dINy+gWmR4Q
u4nH+xHMwKSSLJg3mU6zCFcQfCWAQmnNQUCNpNscZqGGJLqkFjS7jDs2UKXoxk6ap+PPdeEP0b+W
UOP2yDoXrQmEKtwQb2vzHYlvYVcGDfyaWkqlmV4ypteMDs3m55nuRyrtPkAC+cfumc+xMX8EazfB
y+sT3vhq0+7gDrqXL0ybzFWpiiRDJ0cOFIbEeL/DQGYv2dUDw1d//ATJhLaMFx4sYlf3MK9NUvlu
c5aWLgHNORQ4RwPWk9H2jP2W+bTSdLiTF8BHwxqida73FK+pAUzyjOwYA3/r+/gVrAmtcu5R5A7C
ysyhpr9BhCDOev+c0LPKvxVplwAN6UOiRggObX9aedV0AWEKgGoLfrokhjIAKQPOJnRF5CjW7FK3
w22qjYRPbNKo19rFQEM9BYn92iv2+XaYfK8Xq003TIoPxarZQ2rB/DWWk+miJzrJ8idFEGtMF4E5
5uzDI8LIKw9XCJqfJon90vWqIxTlZms7dwZJdpv7ljnrVKGN4MYWyiWSdbQWgkADXGtTSuyLTWI7
9yHQKd8VqRs8+frfEW7qfL6y7VJx+v6NIbDqyCchLb9GKLaZB7IB405Jyi686pGMwcqzjLm1TDZp
Wfswa923CC53+smSyIsF7u5hCSab0pRtib7YRZRTjMrWFuAwanPwfTL1kjrO9xOSOx8wY6vt31Zu
zQftX8pMoy6u51c5/wxZmf6lM336/Ub+Xl/gV+qbamXdWbzVORIcHt8uQkvnQmIeHh0rrOT0tBzO
N3j3KPXTSffDGMYne/g7WfwFZET8iQGQiT7SoDAEOMR3BVDmetw/9nzhgjoqhojX/MVJwDQpZqE0
tB2HcH1ozAXfKZWrk+TQz4XBRAZTAzDmIBzHc3JZNt8GA9N2PY6hq4NoARcF/coDjX/1zLugUlpG
kKoseOmDCrWHTDX2R2LtouG4w+DKmkJ380Jl6CYT1w2Bss3JIRIu9E2GdGxDlqQXik7WBDB7JDz4
So7eYX+nbO9ZaQ0D+EdRIJ8B7EuNrrYB5rVTIWKVNL9pml1gxhqsxaEpPb0OU1QQl/NUdJ8gLFgx
g5TcVDS/f4ibMZKPMMTqs/oMwMibsKOnjBLF6Y7KJWAPBau3rre7vuazw9XOTYnBIYhgszMx1GkP
rmWlvDd2nOz7k9+qVsdkiV+Us2TiMrWof77vTfSYwW6/YtpcRSm0x4ah18B0JVUn0wF8xEtSx3uU
4CKokaB2rjL0/y+DXeGKLk2ogMEkLAUESUx/uYzrI2re1nLCD7PQKhhAU6JM74nhRn/Zx62HFq16
sk5TTUrMv9oRgGV7NKY7ZCxH4bLPqQJIKqhWgupJrY+fheq6tuhF8wUtOqbauGp+cxI2QmE3Evgp
qMkJuE98eYwNdTf8g1LIo7PKkD5c2VgsoVp9UB9a0Y1nT0KKoa6yY7fnNa/+ux85A8ixvnvn9tm0
zqVgoLMr83zkSSLLMrV7WJxYvnOmo5JHthOymYf80WDJPeWhDrL2dKWYZVFvohKzQbD0J2u7PyPn
38VXdcDVmfEJ1a8OMGodWOTW+K9PWVvKoYlL/3UEZXykA27J1NNxg9QckXpuvVuRB2oRhxUVzRQy
DuUrGcN5R0rQXHfpoLvNCj44MoSttr1BsXDU6BbhSFrwSQxbcbprlwW+XHo9C5Ed2mRqY9Ut+VY8
vIej5P+qxQALzMDm8piUdypNjiF2qodNKXCpqZ+s1THqOnuR44PWlPwT2uiOEsY0vEPU2WedTZ+b
Ej+7RGMdNIZnk+xUlcr92f8XXK4FS7DwQA3nmAp9HK2Z1wJcQq5UBIfiRrwl0NUOfHqMxK3UwJ+x
pVri8vTIsmL7utSlE+Y/OtdH3hp34FdesU1vmliBvs00bg+Qj1CW7YVGFlXfugfPVKM9C38vi9ms
DWA2OeOEP+dK1Hcc0ro1xDbwUMVkEAmE+B65M6M/rO8J6hRLsyygIbJ7PcGvBs30+iv8C2xk0Tkp
cYPL41xdYZxDzaLiGzdjZGWCYA1ZXL+xoDO9aGVJfFYWN0gjjlO8cbSZOJp1BldzrWtRsCSYTRuo
jvobZOOFlRsY5CzlFbJSgtSWgidbZiMUOpowySryg1IjF+aS6Uozkr6SvNXHfhn9KLphfd+RHNx2
PV1jLaHN0mC21jjhszxlzWHTUDTizfYKdm95HIDoc3ggemog+oLvbaIXVY5c07lQKNGeN82uQqz9
J32wLv9wibHOkF7TPuFTgBbn5WRzF5kZvjlSEQ0V3mWrWIyU8D50/uc0TdABekSdPy0GnyQVPJv5
tq7Ig01VJNXjzqugSOwRRsX4brgU8oUZ6HhIrZZeCA9G3mMR32hKt+2lX6HhV6tcb+tl+G/LpeSl
oy9h7it3MOmf1Z5o2q9YW9QTfT/gHvFRltjidwoD3Cjou22JNuAkoT0MGSAy3uZ777RBEOVVYRoQ
KYAljkaAH1OT+plsQJpXG9/XqyRYWAF457LCZzRhcln6pjzWcNcUopE9uWcbFzXkEv9PkjfR8CA1
kOuRdTGUtYPi3cnZzvjwcaDN49d3ZXH/00eI0QYntioINrRPeWgaiCDdz4tl5lcfMFSEmhT1y46w
XXrGpVNfmcZcXVLl/pvPtfeKZ8k82iyTlRV/RAdU1cDsGFkoG5fwG8ph3zOSYueUszYTnC3PvbJA
WA/LRgmRtY7ziJwR4khr7zdLPJIuy32VePTvj8t5eQdkNzJKv034dKLncbL/rE8jwgrQkl3iz7It
Qt0XcmxU9p9qj7iAwfs7VSwKnRIGJVKl4R8hwXomHwZq/iCekxUVLZMZ4JlSB6jCQljrHK2arzlx
0UfcIjVq9Jp7m6jhKldjOmbHTXucH+X67X7b74bq9RLh0vGEmFHiBAychT2/OoseD4bzccY0ety/
pzDBifKuWnsQfzU5dwv39oos7HNdG1iwLukn62qdIQy4Coa1QbZEqli3MnICopPR02rocTUcKXKN
fTVpNDeRzmxYs/Spe77mr/0GjJL3CzV0DYVAW41u7Zdk8AzO8qqWhYzQpJBFithlVODlSvVmhRux
VzWywd2/p33i4xquRufNDTQAMLEnIsPPBUBEydCm0gBZHqh3vTlsY516Kz5uWC2CVACkJPx/574j
HhtIN1rx4G35AJqoIFUnFsej3jeAnkLZ9kIwEhG/l+fM1/hd3V9xjA9Xxrx2oll1Ky/7hVqGCMcS
Qbrt4FrXgUX0dAKgxhcWZ4TlR6HwdZWthfnn7jyRbhpPklxEKGXL1RB9weEEEMVmydxA/MeCJJ90
QmQ7ZbTdDO3oW7EM5K4h8hyv8xFmWde74rL46qqj5KgM6kLmbGGbd0T1RBJyGH25zTiEVrgu6CTG
7jL7xhYcg7CSu0WWMjMpwTYkVU08P+Z28hNdaw0ZGUUbHH9sgZzDRmUIZMs+6bwhzOdPGB2NwoR5
nHwRpsuOnLoTrMpf2aZ413EMKM4aX3H0hQlsob7iu8AzFEvJOa13Q7NTLCoQRnnKX49wWWwssp5A
8170mN8+qzGiHfSs129yOFKKqfA6Z5LJdsVoYhJTW/hAjK4cImrdqMybAxwpNXR+19fdm2suxzHQ
qRMWGuq63x/xdojOTWZv0jQp9zWe9V5uBqgVp+JT4HO5z5iiRALAdm0OV/Bt49NtgOtDb5r+nCo8
+F4a0dXix390y9gyP+zMgM9K4JZFJLQaauTwJ0PiFMjYRTk/PV+X6NQAhlsa4XvE15T14qLupZrQ
ehXcfBEJjdzKFqxk4F40py9cdeVG02kAb3ofomYLugQN6CvonMhMKB5QnD79f9g5DHgoKJ9/8kNl
xsdw4Ii61Gb2F6P7dStjPLcr3CvEtkt1Fc7d27+d9N5mZ8BnWppqdjNVpZtt3Nrc55K0zIszY7wz
Kr0l4h0VWKIVOcRNY9vVcJIA1CTHnqSa34phgvgdkNFbkih33pgXJWxORSdGI2cwr3vMM1o9+KgW
A5QDpd6H3ZzKb0oyS7gzIQ5vMs0eHGE8HWpUeOHDxIfzjFKlaWwdOBSyyTuqvKd4QCqFa6gxve9H
erQnX2RPg1RXqus9o9GIDMEtdnOIPBcv4H7Mu2dQ3yEgD8aF/0UWg+rNiP/QylEFhbW2021O9VSX
U7HVJAWXgdccmV3KZIFvXXtMoMp8wmCcjGfdG66oT44v2HXgDDC6UHEpGMiYdkfbOq3HxcHLT8Ko
sliSkoyygKcLRhpnRfa/INFvpOIj8ZZPtgaeEZZYpUAB5tPlQpMcZ84ZUs0biCobNwg/DCcYlH1b
IrO5cH+qph7pOVcPNVEILXy64RU2nQOV03itjZx8APEskaflZJ5rSa04AUFqWhTI7BlZpuJSMoDT
L9WtH4kw2wiK937+2ihvDABeIcVlJ478zr6ssx+HkCM2IF59NeIWrIAa0pfYG/5R/NjhRBQh3+DZ
E/28pRZD/gz+cnbRiF/BNjxXnV8rNa6tEqTAJkqc+kKEZOJW9ghhDa/ok8QL/ce2Dh6DiEZQ22Ul
DUpYm55JbKO9TGZZOWTQ/1rYJMZe9VRIMfJ5qery5nSFNd1TtGgaCJ5kFfrmJo0YYvO06GmT5I2R
H+hGFdDFUgW8STOACFipnTpjDDz6ZEpqYIDeznHwLGEQc4vymJ4UtuNrgY6XfaXletW6Ui7AsEvA
EwLLA89IQKWnsR7JWfBysQACoRxLBoDLSju78VI/D7wRgRVzXRNhvwWk8X+OLruEs9lsiuGlwUJY
vXACn3iwLy7va+BIc2pwskVFXPQ3gCHOmPBE2t8dsVlFpLa3igwM9iu2O8GJvx0rzieMuB/LytCH
1dONekLN7Y1YiwRv+oKGjgYPXVE4K2ncEK/PE09jMfQfeuR5QmKgVZtIz0fuWz2NtiUxezxAo/l0
zCujwVsuc/HPH2yvLC1+/a1TIEv8tXbYUggHBk5m03F/vMhwLSsqrgK/Kj6chCKWdjeCHgaWcDEo
SH1fZwu5rZ/S3S+ko8d403TEFl0SRs8d7MWofWpt0toK+ygL12eoD+3DtaO3cb12Gq06zggKiXi6
laYRrXTFuiCJIXs08qKEebTCT1Cn98M9yTqm7dQshjj+UDRhDvvZW1NpaoMTZ76/XzE+S8hQcFZT
ZSS801qfkbkQloC95LwwpmehHmPfDufEN+AwnEtIROgVD1b3UxpGrlxsQpV9Yd9++uI5Chr+OvPO
pERg4DvvFhY5oEnWnautUABFNcfGTmrpRHY/MdqgsMQsiPqzz7xVvvRkrEmsDWvQziT6UGSQ/xgo
lzz6DQBKqRiWnNbDPNpPhF1iENQ4lQZD79XNv5v9D9f2ugsX36yYZO3WrLkCOOlHju6dO95vnvXf
QyFg+ISnEWu3TVRdJkZ2VWPvXtQzUsh6Y5wAc0CQHreY+VltXsnAvXFmnOthfBpW5uKyHNCRMKEN
hq2Hn1KOin9hc44rl4P26rWJuuYpVXPNTIsHdFY11wbbSAAxV5kdeJtksvHCa5Udfo+E2VaP8Ot0
HxjeLwiqWHP86DI9Gn7zDD4CyuonFe7o1j+ihcKfqwh/VIfq9TKpZ2nEn0WwOhT6HtdKn1oiT7Ql
mKhtDR0umOQf9KkfxsooFTpSRhtPsb42Tkj8PORuDBBdQqm3FadZov3O2HNlP9WnFhaDikUadwWy
6wuiBmwVh3DZjTB9vYwLiWVpXQSIoFWjOeJ24Z2g+V6UZdg8wLRXPsueLSkoQVEcEljiR6rUmN+h
94jWj5j06tx9j76n6DMWHndAiSIp3hcOjCbIwVuRICtwcYMkIIbE5SW7WOPSp+CT8rCcb0bSt5/f
AtQLvY/aQnHWhwOrn3UHzko0VFmgKFewqSgXmgWreIGnhDdhTtRUr6L53HdcCAYbfOLKSPaGEcd0
gWcjkB7/nk1kCq1Pm4YnLIWMzjPZHAxzwhuakUBQ4WD/8MZUIqT8S78lwofC/YdWeKKSrCbH+Bas
P2YHDso0ZgmsKrkf0eNcjQ4vCj6oG/eEJufmbQRWj98iYL98EuBuJDV+EyGWHT/fpXntag+OL/Tv
eMl5/7QOHNU6QCB2L9NsT7kis0aarY37mq9RC59dh6lUSbnXZb4doLmIQHWoflZ5VWf/AA6WIFP+
UoWJ6Y+lhpHcK8/iQAkyuSZW+m77/+20G99JM4nyeV/erSQPOVdDVpBL1kSq2TymTMRiciJW67f7
c28LISzh+BG8oU6QcPTddD6GWS2UbhXyyIqKvkfDjrAzDhCNzFBktqFWTLItZq7bI/DdjCu5Q+rg
zkf18g+ORWI8YqEz/tiIZ9SPztcuFAD4Xa+uxjkChFh7Rrx6moT72JmD1CzGESxVe36TDX8vhNix
hj1DfbDaNXZIG38nR4Tk/UKO9hdU8WYB0LjGRqja9mLIDBFlXfYR+yWPGxrMBD6+g4sw8QnQQ96I
yrvS/jxp7Z7Bi0NwqCvHnuWsyCSZerba/lhlhoVvMLIVsgO3BZZ8/IU60H1hb+37YBvzREIqRWHh
fzupFmu73cvIDkKtbXwguTj6jsGGmOqQXoHh/y2Mu8amEz4LZcGtPGmNunhq3xOeYYtJpAPWfKHb
v5xWsE3mWVwSQ8BUxAAl9ROIs7ul7RfSnq5CT2Kf4rS5eMFqb9Un10hoccen307sgCNJ1lwfm4pu
oaXah0PxE6b9V4/xDol8DZz5phkB0ku/RH5Q3lO4VoPnPqEZjwaArp6yu7WIZ+R3oALFJj5sVhFM
MJSOzr6lepVTK3jnril66e+tSZ0vPDOLGVDCWLY27yfCrNioxEYn5SJoDiur8O01Hf0ynYR076GN
i/ZJCcdyHekVSwhazWpwnPVyvJIPcmfpivxWa7DL3EHIfb9ZUdC5CsSU7MTeWm0CnR+Mg3G7Q/6a
9OEDHdzjOCOoYGeQIhcnnxUGIWgAohwcuR/tSQUEkpheZXhrnieibIgToVw2/01Ltyu/sxTPD0c/
wJbFmp59EWOj0xrp85s15EytlUZe7xVEmDSPP22p2HXbXGcO/K8xpl6z8zpURE/mQ95RiajotcIa
JhU05jdUy5Ylc74Su0YQJe2HMmPqVcd0gavl3qFpN3m2HMbHQFfxVAgr1No24brJccfQyE8JhmKY
wK5fca8DPDXOET5BNee9g39lJrowX69tdTcAX8D77NERy6bmjrKw14qB287BRC8kjfCyTO6X0e9g
T8z9E6pjybDddJmybVY3wLz6d4WTvBBjKiImnLjPqQrDPTkbeKXm7T8uFNhuSjSHxx0yMOxgGbrN
wTw3Co0BTTDH0eVDfL4S4La+pD0tlK3nnVfvnhO1xvY8U4Dqmb4xwFi3JMperZoxGF/EfYKACxjv
2cJSoNz4GGShXX0DJ8ZRvSlypeGBfDlaJgtaQqChqOdXdZFAHXAAEThp6pag9h4DsS0qM9vRUW9v
uE3ITKqjdmyoIXhPHyUfUxjMce81AtDKVF/WedVjsGv40SVVIJQmS6izQRniEVZLubQEBX4S3keE
hXxKAeH9vUKEIk9F6ZxwZZosCGdy5J8xQySWBDHS57Co5u8GuxXcN0jJ0Mea3zjt/HG369TAn2Fp
9MuO5OG+pAy28mrTIHVZ7+RiDYQ2pexoPhKBKNI5tRxkcwTSv+VvgbFIhjxKWMv0T29bXIy/A0TN
6vZfHTQDUdKoqIdtQFBwloVU7ZlwTEq4YYqB9oUN+pt27Er7LOgbTV5wDk15++jKxtQq36ANwiu3
MLlNRnslJu8MSWq3THrUtUV53MNnFN83TYqwLU5wFGEqb9L1Eb+3IzN95BZnDPHQbXnz1PS4BKpk
piWFoZvprPC9B4IDBusTcpagjmNBwqAXq8Ow0k7xROWmZ9SqJCTl8y2JrKFy91ZusjdT77WrYdTD
szFL5ww+VBoGso4+d2PqVK7+GKHgo049mEg5S7zMlVaQTt9iLmEUZrVzMMW0jSvmDnkii0KTc0ZW
MydFhlozsJmWGhQQJI05lsYH9TpSj1S9McJWLHTAPXgDxmxE53KrSj4nzj/E19RnwX7/Pg1rjGe0
fbv3P6d39nijCdW11L6ICJ/+wT+yERQHkTFWVjfJ38rmTQAdw2eGL01MsjK3Dx9Oo9XNbfZ3hXvU
oWCEcNXL5QUfNvdmbaHWmUnoX4mKiFhVrYboy+b5q8ytOh7uNXgMrAEaxcr4fqqdKW0RT2B4F7H7
qkDBsiC5XLlH/HolJmT4k3ZnRdafWYMGv4vlqpn/4ta3cf0UXahF52NDO2Di1FA1G84G5OgxY8R+
nJyrEveb1J9KPd4Apb6FqZCwN6lhThFRyC/iWa8sZ35IUWCQWnEttZX36cHkCwCM5StOczkkBISe
BdrvbxPVRe8ija+K11A63VUgh7/tVTlCXO7uJYTCxpBCksXWQgkosjP7Yk2WSW3HhZo+b2HrsQA/
SRsbZ6vJx7ryXsqcYhJQ3ei/6ThnapIr6Bl0hlWQYZD7pwUL09xuyl4Ika3ptsJGK1auJe+E0SEz
aCG/G2fBpQxC7CT8mKzpEHcmEX9N8HEwZR7h2VUcYJIp5mNVlsJv8VHqR+pXl66qBsrR94eKpa5N
ge3t4qoQSFC1MnYJ7pojm6FL+j0+osY3jPRMF+ed8MGAxXZGz9AQPRu7lSM/UNP6vY42B7vj/MIH
4bxGdq+3Rs3EBBsT+w630nmwhIHAHuPzieV4BE1/nEEiAybemINIXDUJ8n57fPp0DCxoCSkn3uQZ
PGwdojPvcUqQ3xHe4wKzw8pClcp7BQtQP3DcTQFefFDHBnZ0+6awgSAp7nZ4/+iywaB9cQC1xAfY
5gkNTHfpmUUPgD58WfOmbCjBB7nDIJ3j/R7KyQrECTQinm6wsYiporbFi1POiW5VuQQRU0ezZdRG
8bknuY4bgkA/16jMDeShjUP2EMuS+YwIhcRMRQP+OQj82b43kytoNqbFQmqiFW2aIJ3YABwn+dw0
8eCfFv6q00aPVq9vNJluGYTprZ49WGQVHi1SjswLgwCjdLqectuu1JRdp+VLVT5YTaHg27RwOjBW
MoawglIGCz9GLICEVWwZ/U0gZKOS9Kb/lyVNm6Z2UUVRMSIdLgQTsqLQvRh9lMJ6Lq46o0iFYIzF
5C/Nb/BQlpohZf0zk9+TMx+ccWXYd1mXN+7L8LiXcx+zvaU2G8J5Vii17VJsB1GIOdsFtlXsmQsQ
R77PCZv5ycVRtETt0RRn3oTOJd+FRq69z4LIq9UcYdDRI26QX1AH7Pwn6bkZ6Fn2lxSjqFzbzj6g
sANU/Ak1l41JyAxKldJPWohW0QRyYHYBW+xPCqkKRoCttHBRz9uznQ7J6wQ3Y4u/OigqMwyA1uyj
tQxMgd7ykbJAesm57Y+nQ0qIpkx5XJKZTQuHXC9uaQix8bwMkyqwGykfCLv4QpAewhj85jJeaDlq
C+BmTyIkhUeLMK2hON5lRJMjxiMYvLJRoP3o5foDswpy57SKnlCTMM9IuDlP3exWHfDO2+H48Mjo
CsMpZfdqd5PIFwQOYAXDMoQW/whWrTAH4K95h9iu6y9wzmeQ8yXXshvvQfjFULcuzOTbwLpe9gAo
IiQem+1PgqLsb1k1F8TfwgkJ+W18cI1JtRAwFR1Lo9FK4aTaxM0ilKUUYYtox00yGKI3+GnWgV1R
8TC8Y+Cn86Ecz6IbO8nAXh0PZw32ATyxUQZcnfQZMgs8YTIaDmYD/do9/OaOrf1sYuef3aBaH5/T
CL+9k1SGg7+qqt4lR3yDUH0T5Wep0tebabA6nu+DG77/Oy9if0OZfVxxz4lJXF98slMGqVap+N9D
fhIQF0p3fubzjnjlINqfzXTo6ZJ8l69gtsZ75jp38RUpxbRmERV/GEvFTEmsU1kkJQONE8UP6wNT
MKvypSiquLXoj8cZxlVKCEm1X9V4oCRZ7xymUFfssv21TpStITRdGpZYHxiT+UJcm3ez8LTmk0a0
GLWyTydzIz5M3n4OjvuHURkiZOPdtfr++Y/yj+t5myAeH1otzkbnvdyRI4fuE1lWJdm51HEPs946
gMfu4tGoPrRvnPv3OHHjtOCWQCxZRO+K9sSYg14pUoT/o0kGxWtp5JtQtw4MrhecPIxhyHLI4UCg
cFq7OIyLb+avRFKThIbZjs3zVnDck4z+b96JYdmF2dUOBzGdVLHyPeyA2V378LY36Z3rbJUgl4eV
0caZv9S5Ax3k15ShaxRfSfRnLt4hyMydHmxfAtlktMsHWv+cpUB/HC/EikB/Ej5ZFZBpufmhCPlg
Fpr/j8/TdrQwHMG/8k6qBOM2uC16Dt6iS4s/+lQ1gbpYNSNbUCY2YJL2DhYeM7d10B1iBT3+7dlO
J7g5XSw65k0PBD5fHEJHANXeMpE/N1EqoRauue60pJh693mehwPkPFCW6QT+6BzY990R/VJJ4FRy
3GYj3vbO0EuhpZ98f0XnbZ4aIPcMCPpvQmo3o0SN4VLD2odJsnzzc1EPzmCLfiuaZrasHLAZYZkM
FFr/RHfTOPInr34nSEVIkiNNEaYa8wVGcCJ1WkLYh3YU/hahk3eS1vObFOKNri1KpyHa+PRpUK51
SgxuPXrZd0tioznxBYzFRC+4qh7CN7kT3gIgH0DB90IocJ1xf00+nNGOeteE8YxxgXNOEhvVsT4q
/+ESUbdxhtiF3K4alxQ3kL4+HTC2MgqeFtfcR+G3CnHD/nYZkwmZRMEd5St9CULamkoXwLHUdOIm
QAkObEnwjLVXPNNgs06RaK+BV/g3nwYxmUlwUeaNSFX7W89z0AqrLYfJRDmNca71fkTu59bZGp+Y
v13A5qUwAX3BUgEE6nNrriAyeZCogHerVDDrU+XAkbjdTqCje6gUciGfN2oy+YaanUKS0ZP2XfbJ
ccLtudETs8bvQmB6AKZXY6kIPAbzx3L/7SsZsneqwnc2VVU5h737WzpJkfnZptOSWKrCc4Phluy9
jOocbsuL45I3pd7CW2cHYTXvlqDi0SUmaeNM0fejmsfCuzV+J76z+WyrdJBL5oMW+Qlc+SAuzvHr
if2Xe4ZokOoTYrav9FRVpunE2kwg08mdXLqHL7aYsPVsXiPwTDyPG5M1YCPQ9oSLy8uEXvt6yOFM
///Von6B60nFED2+zfljLFiHhD6a4EI9QNL/G4VeNgva3Fs3s7uqifyOziZdiBFEbsu0vGx1wGN7
C9YxEt0UStIvyZH5cDDzvtRI1MNi8QIiD7Atq3ib7rLFibiSzLP8Wh8kCELLlIt3P9jtKi8a4y2z
3IlFZPUl+ssRzJG4yp1c7OZfb5I0pXjnFvlNg9lWOWcSKn6ZsbUgd1Fg8yTZ699huJMnLstx0pSl
an+uc94+qh4J+aFIzm8674LZA3ioBhHLEEC9Baa7IkKSTdVHdt62hKS5soTEVHxj+wlxDSRwj5Kf
O1RH6LYlK52jAbMlLzQ/eOBXSpHQE27D9a2AxA+Sqmmk1NwwPTxTgd1RI+J6DyjB4Wwpba2uwClg
+ktLchPpBh1sKqov/hTuW7EagCEgEcwJ4MpbuG4xrIZ0SqZcWbaULVIkMaPrTl+i5z5OMhPcW4dN
u7ujF0cbFZDqNSICnIZ8kf1a1rjxxbDOrsw2BkUFszse9gFtHfTvVNv1B7jmDvNKeuznIBFVMEYD
25elSigSD9NTNWl4taRnn/95CwEvldJHuk0XQlyZVL4MrLZHJlBwLdNcF2AAj1jxhpQHIoA7NABS
Ys/y1wsH6H7s7HHaSMX+NN7gRXdOF2SfR9L3CzkhkyTPJQ7yukzEUSehwRfOE+mhP1g5oQB/IjMp
TxpWl2SUSiCEd8efqLBE92+yLrQEnyAjv5/Ih7lsGIp0Vn2qfd+kRPFd3jeg1etOcXR7elgrOU0g
tYno6/bD0EbNgBhnktgV74YsHQnjXxxh+S+rKU94rzkREp2xXDWiwdhmHHuKr41EuL0CliAPfNVX
gZ5iYmoFS/pqaqr+goD+GH7+r/h95Ue1lSCJO2hwR92NQXf9hJ8tK94N3qDKsY+pFmQ3GxqO1Dyf
tHqP3xTR+3cFOqhzjO/LT4cEnfc4AW2XqKKjUfCBMy37TnwodUVRhmf/ZE2PMGL09dokx3xne22J
+nwJnu5zwi2Bwe+NCw5KknwXbJI/6vg6I97AU9jZeqVfqXIVIzZk9zVF+Lnzd1iw8V+spizcVg6I
I6Y5eCjfzbdNTQauuO0XbBhxMmQIaT6pAWL1DfywJSI6NqNoRUKXX4iUVU8JLd1atm2CD2QzeE0F
DlhT7QzFOGN2L3EylFnPHKM9nDbh5SexUwtUPIkAVtwZEpnKDulqU47NRO4ORBJJ1+j2RFVjQ+XT
x2Gp8QeE2VCFt1R0rUTp8qcDoP20Wf1Z8jA47Icdvzy/o2xVdccZbKehmTDDzxiW2IVxImFzKa9O
sdIwjlqGRxKjRWawjHqjpbPatXQWhRmPwd8EgeRqAVaSCZDN7OHskFgFZihaVMrhTUDkHP0qJEiL
g2REJrzO7XxZirXKfot/lt4naFVCcHTqORp1m7vGk+YQMAXumNLivvLp9hf5sVnuMZLAD7awfvpM
TowSipDMNUs3bbdIazEPGptwPA5AUmikEB7/NK/m50fZ/kvUpQUh/BudyAOwzgXTgb79wpYwBR6D
RE52IsYuefJphVku5Vhw8S98deAn7d1+j2Z87Lq3ppaF959MGYAB3GvHtqwE/zb0SD2bHYo9TzEP
iHxjdvkJFSuBPRN1Tfl4e3cXiONvfTX+oDPVcyVpg8PEIvpoSUTXPrbqo7xxvfCR467S+L3sz+CQ
uitunZShqnBhIbSzIPIj1iZD2uXfeCyFH/WSt5iJ09HQ78NZuSBnKauvnGPfWbOKsaxhzO+neoho
fmnrb8lOBLRNZbM0OIyX2oRK6SlcV+qbksbxwWP12/e0tMH+x/oskxbdAe6l2wo2fMMze7kn3o9f
gvwqhAus2mOyu2yso3MoMl3q1WT+uMIDNX8WloR3Fa1remvc+w/hv2nAltLwC5jewLtGKjeCpZHp
iULZFFjMyXjinCmZE0Lmoe++wqKoxD8YEBjB6ApHrHR4DzE9jbTWGIcrC4xCazDPiUUP2KIW5sV7
cEd9qz15aUKj9WMb92LbPUvIzg6Obxicn/6n5eW5wavGOkHgnAoYlpw2xpKLtr/RoXxC785NxaYl
lxmcy85oba5ZGz3G86KFTgRFj96fMqDvd5clnHk8rqyBo5Eu7yvxldrAmfOApvpc272VASsA8tXL
1Tiqn7nWpAP1lP/0O8Gr0QbnA46rBNWqbsVoJDzZBn43+jwliBj/ZCu7350xZeboO1mF/3w6Ov36
KQi87u6aee5Qdyvz7qVqi1GMuERRP3fMFdDhraYhneluJGtr3v2VBfi0N3npL9T3bqfRk5QiUxK/
2zdkPtXIfgyNB3gLSeqkGjbdr0H47HlxNiaO9lz9FKgLLqD+iD1UG0eWJDYS80bejU+GGDKoOIXl
KFAuOp7J+jxQTAXDt0cYySbTxMW2GHSJhuNvVG1a8J7eGQi9eaijEGaEE4KvV9wURra8CS2MHk+0
Q3K9DPqUZ2SA6o9pR2xOSDKdZcZj8zO3mBrEDWNyQFhvE1m56kwSKAUgz8OEQCcXzqm8c0ASXcqj
9Vz7/vyVAM+Sbf1L1WLQgXbgU+MBBE5Eb9HyrJCAFl1Nfz7oaRXzyWwwf5tmCyYLsYrO25MQh0Wz
BqBqNv5HGIqCmb++W1I878l3Lbw/v9B7yXrxeYcEIFR+/IJa1E+AGzAToYjRE4fJO+v4TgKrFgY/
nC3um7TnrdnWuf+Z4+wnLTEC2XnKS4vnDH0mQEC9+HzWnxOxrTLqbqOEqgmgT9jkpG+lTzSfmoRo
Lv+HUhUnpMjDcAvv6QnGPHDtotfp7oVl1mDhFO9q4xauDcSMsiuXeE8HEnLjl4dn6Slm09jGq0Of
DwrTmbWcbb1/uCK2Xqlyo4bb79AWf5TUBZngXUhFZxU/kjNWbVolFeC68ngLb7cETzmyYikbXZ7M
Y3Qpn/ADYGSKoesSfspC9g+Y9DBHiMlajvYGkTiSf6U6WEPupOY/3CJKqnlEwY24UgtGzdygHetU
AgR1nkk6pfMM3Kptx36/Ww0rzxSIgel+J0zGzp3oNhZF+pkDJ9S45BXNgv02b8LXgRwt/x10ijOz
B50VhbYcJIglle+tiXAiePkqIOjwkrc3O9kwIFTO33roCOIF++KrkM+Lf6cZDzuuY3+BeW3e0TzC
7VACns9fm2btWVGnbQ6i6BvcqE3eSmQN9moqdhReg3XUv29/+3ExG6SK52JrUU9FRSwvfb2RnfOC
RuarjuMbGlER8YAyEc4JAVmCUtpCChmL3nWV9H5QupUMi8+iScnGY3wDGfG4Q6BRiU72slqGPWAG
jr/zmF5iE/EnAqaRERlCHoYakWn+4gnL31mD+42L5ka1zH5TSvH8w2y9tH7QuMXpkMWOvyN+MsNa
tUfbQ4Vm33dNQaodG9Qjxp/iTeNacrVzGZ4L11p4kl+7JJIA3jae1XFn2Q0YK+78JNovOg19hsVq
En1VkGCQrvc3ppnKOZxrEBjcLtR/zg2KdYXkTNPrvXTqOPeDV/jaBKoNNLHA9DMB/KRnMMp/vHqE
OmlS2Er6SVn6+qN0+Ivdj2quLeVO+M51x25aB1Wg/m32/PMUbFAWXpiqFklBX+wMtVZ82TWUwVIi
pAxqk/W4scuLyUs68QyMpwwjTPfsfpeBsQC81Exrc1CjGN43XNGu1QpNYeH53IVcMRmBEVnUWObb
BDQd8B0yLfGnlWfaVMUUnBy0+SBj0pjBZkrCWn5t4ASqMC04ktnXYQqc2pnm36JShTveushozETk
dRtBMi+KqCqL+Yn/3GFS/KYU5J0/kRDHr2FJ8Hqi7RT/Q+WZIFai41YXlrOyZlOqkNACMUbbofQT
zO1LUnAynIGFAkQUM5X5jdjYBD4nGIwxGGLj2Gks4JLos8DUaMe8fLCpAbLsF39iur8nfzfHoUKY
3UxviXxA94EibSm9KtCI4rDIZUmHPmuyxqe/tDJGc4Uw+mTuwOhErzcdaMUAloA9aaH67xAdR39v
1HB05Np8z3ZKGxrzjuyryZsJCU0Q5sh5YhTunt6CLrqyPIyo9n/MD0AHAKviL0xCL/RLScv/W3YF
mVVorgcqWH+lEh/VYzU1s5/hg5/pNzvtuHqa/IhhLFgZy0H5BATnhPKp7aoCFLLQqqO0Lgirdfty
oWKeskmIlZaIvRdBo+W5xC9W0pENtp0h67pq+jasAMOp2lPv+uMs8tmK2kJdFA8eSMUmcHKRtl+2
sthQq4KLKGcmwJFqADYZoXh5JncKT2VcQUGImpJtJhT5Nn6D5Pp5cb6zegSVOc4hBck/0QILeK6F
CBXzZA/g5ej/WG6vyP7E5RkLct0fzZGUqYfvBXy+U18gwa1VP/JD9xea6DT8IJhanlZsf2N1rypw
HHR37SxHXqd3OkVVdyJRSxZqOQ3ytRuyYr8XtkxcL8npni8xT/a3c+Fr3G6n75On5ez9OZ500LZg
c5HZ671QZ4xPUTV2NqwQcuF8mJ4ArVZPAu3VjV8xRtNQ5zlVtIMofPZLGPNC5Pdo12i7jRtkfKRG
uhiXmm61+QkvhqyvedNe7plbbqV+4tTdhL4/6YynvO/g6H+fd2bFwsenu6BCib3dgMEFSe1HauwY
uanDiamtfauflEB5tjPR1F3jy1aLGNrxaSrSyHhaKQHek2r5vo116tqM6AQT0XM+9Kr7SsraCJGH
p2EikH3UoAoq0YQlnUNHm26ors7A8jGwP6onFX4QoD4K2r8LLlKvG8sSkCJlLm/gHDIOkD7MI29j
Fx4EiiFKqK3LpCas5i/pdMVYLmU4Z7N7zkUxpz8VaCQTzn3rq1MrU2zrY+T/vo0yaG0ghTJNJCLm
N+vzzTq0j50zTC4sT6HEjQnKQsg0dsYHr8RBRiAuC3WclSgUXs4kuZnllR2maD+kymLKgnF1whmc
RdfsY5j2Vpgei26VS6RNnTv8H+l3yzv+NCRsvUn7sSAnpYLLXNqQ27ZUFGv/zSZZuquIzEXTAt1C
XPrmKXmuR4Xi+LhC1ZfRKVPvDWqucewSWYHHn4gbZtpra5KqmsQTo9PuLj9ZbhpxefEshheh/bbr
HJjao4SpE3fPj3d4SYfskbuhDKT2L6zly7hoj5PbIB1rvuAvvkRO6dQFSJMda4fLq+vbH/N1xHoX
by2iwVR9Q9RPnx8cmFhZTUZ2bT8SNpiwHHtCwIzUn72X+kZvK/dBKqtaTFtqajvG7pSSlhn0nii5
UtDfkoBRTagMY2MbkUR09XniOC7914l4s1vJ65U2oilpRhFsI2KRrki9t2C+keAbSQEB9tvDhiFh
yV+QZI8zOonwzHSWEY4/h8ron551ByAltnf5pKT5QSoMrWSezfnbBK3k5MAZfv1KcMKe7DWqpZbf
1kS0bhiPQQ7GLK1BzuPq06gEDqpldu+splHfCbM2H7XpXp5MBT3T3Bvm8zP1UVeM4X3HiFr+kXUj
/oby4xSlZ/LNWseTABkKt63ID7fhsndvakfvEV4PQH5GuxEijqDFd4NmLUX1maK2qQK5Kt1sEZPP
DE6v0pNAYltn5ExzuhI75+ytHGJC4fv0qLjONctnIZMqWfzWDlGXuHnXHINl4VL/8UzpS2sGFPCS
u8gIxvTlbKqcPTbZYIqEwCJYenRXXmn9sfsupHiMsh4cLjesZLXYwjwOVDY+czd0Tyzem+LsqmLf
94iAqlp4x7YtSmVw2ea3LMNoZhi283bgAz7+61IpeAGs/+tAjX+BP15rKo0tC2zhXEDYu+G7N2Xj
lQJvoY6EhUwiVeEdFLZwOIcY3nCuY84EK7nCpYFEYRNjdz/H/GjJ14IXAcRRVmE/Xzeg+3p/SdFR
RXMOWud+sz/urdZIeCWFDzruVoNlWsRmjsLyXTqkozWSjaksWNihAaT9Cy67cOz+WaZnfj5b3IcW
LjppQwAQcYbxt3LTDRmHn9ltADyxxU7gl3cjunOq5yn6XnE34VaL5sKcz16UxXXgCJTZwe3mWbYQ
MeUdHmYQWsSmLhndwkKp9mt3zswYEt6KbhJcT08+KVNV+Sh7s9sgdRYfQgfwKuR3OLb47aCYMn7j
GjfjG0WSDVVO3LoRxq5M6WisTL44mIvr2J7BPhuaYhl+RwbCVP/cOtOpO5TysUnGKJ9ag8e/PN8n
Q/+FL4cLJF3eiwRo6zsN0pHW7qMgbxKvo0N9cdKVmtwbnuV6ehXjKnY8ql0Ne2wb+PBPnCVfSjXW
5rU4pZU7D6YgIO/wo2zKe1gEROasBArU8DF7nvezmRhggT+LY6cUNIoXu9CaIh5THh+pvd3m6Zdg
2bhS3l5l0U8Mr5Ug3AbX/hF8lOqrnCPOIff/SOiv5XCxujOX6fh38PwSGLfP55cnqk/jxeJ9tIXl
GwErocu9JY65cyjnp6HNpCAZwVu46FX5QheIcAusGLfTGTVawUsDjvwWRmUMHQBnEyWj8DA+lYcM
kBzC98fRjgtfzxukYgUQuaaqbhj8CqUSOClRZsqxIdk650xLYSP5oddptP5C2XIe46g9n5RuGdOt
lW1cpKlcn6tDVJpHUXLC4V0isIlKmo8qRSzB7W4M753gV8gROixd02eh4Y2DVuNPe3RDQD9EAHH0
zU+Ymg2SBpaTGw9pRtaQn1Y5PFgVrMLzAkzzdm/qZKdrAHFpCYS9CpFrNbOfXPifrshudzS3p8zw
Y9lqmLKkxUkR5dsrkBk9wFqQc4i+Cryg4W03g4yNZkHbbbSV0y7/j5Sl+WKOQutY+tkKLFvt01Ml
FstgEhvKDuLLKS09eQDzLg2LS391maJZiPP/VM298AO+znnaJSj34yD3hOfWrQA288IfvFUAfTuK
8EPMVB051GbN8NJZoD1UvQKIUGLTohfVa4b348T16/fWaY+i+fmZFteP2dAeb/OF+Oz+jcqRi8nW
abkpEMssmAWULukwwcRWKb/sBgz15P/PebwUxebkM5JhB69qA23G8yyTPo4p214Ga/na3KlI5Ldc
e0687D2YtdRtbhXfpOI2WPRDE3HXY0H4st4srZVvATaMI6RCQ0dvmeNoH0xLFLN+JxQI4OZp/1rC
c9povU8XR4J9YIVMHXvKaWB2KEXf3OPkkL24qNf94rbgrPA80kPOGhGvTtDFQZzvXb8DkvPI4kea
6Rz7m16rTPtSSwVh0dUNqjHDnzC2OTx6XbK2GRuD+9dPNdKRfzijmddd9na+vMrRVF9ZlaLXUxwn
I3Acg1gFYexaYfSOcLJtpVCWpFqxsO3ZfuLjiV7dmF9N4h/7UiKajXPrMzpGVV/77jhVOZc4wjDd
ZBv+Oikwys/k5odTmZI7Xh5j/bgtThP++J3vcgLJEROQuhd9235s/xdDtSOS9nf259s/VvUt/8mT
N30bqtGlPMCEGxb14OpPEuZSwsYh+fgVniKlOlTAe+ZsL8wBQdJJllOHoGehAP66bWP+6OAMm4kk
KqSA8nQ0VKY5LFmson1ykhgNgKFIAntaRwNO2x25dGEWKWdBd03yqK9luCP6DZc7vfUHSYfDDQ/l
oovZ1Dz4uK5GL1qTt4fP0VFjR2LpcC1PEwZzcLR8fIoe0mWjmZ80WPXvCowggvN3iac3oltEsJxG
T16bh285L2I+vWmYhDlanR1gPXQVd7Y9h/7qmE2UaQzVZZj4CCOM1Xp+UAM7tJ3fOfM/2/VMA6/E
2/1Soi2EQWgZ6/AVg4Jv1wqUSFwH8a2xvWITTyQu49u5si4P021Bsjj0v8AYgFx2t1tbl/VLm7WQ
80UOTQo6lerkLgNusGVDZeHEDqE5rkYF8fgcEen8hcEnLTbtlNEbnV729QtdrWeOriRXLcnSpjfI
biKwjshtvdn8MimYwsWkLcvCEjyXj62Ay2LWAKYLeY1R9teT7qazMi5H/447Y8nXrkF6LCx0PElQ
Kznscmrs9DtprAqpQq45+ZRaZO00s8FBaxKIDWgSGnqGh958bbPlA3bmXx1X+1C2OCcqBdIFE4fN
vQa4vdScufeuDljM7TZ64U8gTN3MSuVKAZg+eWqxOTBtHbzamPHqZ9XjNcrZ93qNES8HGSbfbim/
xnjyiXCrHazWAVtyjNGrSN3UJ2u0hV5SS7EcaeUFm1k95Bw1IGV352UiwAVZWGuTwCnxQ1n2Y9nv
N76eBbkMQSwPST6SPSPUpdixpovIHvaTnRzS+a3oDs7UlQ01KzE67FNbmsfpJVtFnIxlqXz0Y83B
5EsU1UV/I2CW+tKbSfgwADxXV0yJk3G/dpp5NAj9P7t2U1tGxB2Nyux+x4qjsvbrpHZBgyPONAh1
duwojASuJETfIh45NwuvpJvQCZrhllU10+qKV2bzeKd3Ku4i9WXYOmZmysNL5ue6suAQ4489BKG+
91jfsaQmILZjvLWMqSiIncPPGX277MaBj94wT4a9HMPwhBgAUFX1fQNlnh3SBEklgmdsUebFkq/f
hRghOQcZNdwwPYd99Fxtm+OgNbOYSd39u0YrwIb1orG1r+GVwFgEiukjA+kyhMBg7PWKn82tdzNO
ps/+aBlCfZZXshfj3UlUPTuHmdnR0tpcVYC8YPrQBKzvGmgQf30bzSRAGrnP6pFsgpxVYrZxCPOV
TPjmtMnu9rWyy8uW3tMUtX3EowEvoMZQ6QmuQ+8ND3ON+HBQooOsEcShewNorgimyYGYUbDhDOIx
NROvbZx+spAUp9cpoXCfZZUXz0zZdIhVZmdCDJ+LehqZKSQdraSJ8Gojtpmgea/6bEp6Ds7aihi0
M+4fCc0fddOeggWQT0gnvOXCUkakEZ4do8X7W3pHNYGAlFctBcMSvF1e9NrnPnL5vdq7jTVtyT38
bQvxwA4l8IINfcM0INNJB2uuPmoZrxqh2AeBWByoHsLluwYbQdpWkfLD+dB2hsKkRHmcLVaYvbF1
vn4vr0qDrpnaTvrxtUHhrNLKfSdddY2/ehPw7Sf/nJNa8OcBi0qSIk2php8W7W2mKmUAUuXoN/1u
iQ2LC3+/kLJzjU1z1zLJLn3N19u1JCUzxPDxHZNDDZVvVvuNR/pxJD1y+EN3uYUjVTg44J0yGRQ0
R8OPB12zMfqpH69uAxdGMh1KIAPD5lLmy3/ITFUeVYiDrNP/T/t5r3XhL0l/muC3UJQZraf2bejT
D7CiSWjcEchYzlT4wtkUOJpwGImdrW4j3c+3dcd5UUZDx07OhqscKdiSiQiGpFAMJdCCCXJHUyo4
KtyI/rhwzQxkpHhxmjBJpDAaSi6JzAq4QLUEVeMD1XuCpzCMZUHr94yqte5EdvQkN5m/SnFZDEVb
X/CSt/lbHiPsF1DNI4Jm100d/0/PzDSOpyzlI00ltTyxdrDrzbZOEa9LhoaHlTm7pvB37JQX3GBw
coHvPNCxjorG2/NiqAK620TQttkHOzEX5m+GwQEvyFA2zig8UKtQrojwq6brbsGZ6pZ9YJ4bUAhB
K6w2Y2t6jOoS9m/4DA54ZACJed54jWGRiW36p8AbhSDCGHm4I0c40tR1hRtgVCi/NbSsIVIvqpCL
LMGbxkmr4ipyNpbU5t40+Geq78UPVKGQ9QbNoNyg+uZyOT7cTgRG72Y4eSIzsMjPCV7NR6FRKE62
QQUYRMJtuP7TkcCxqw7VDWVoDSiQTx0bO2dMDSGzD/gYtsY6yfZ4xF2Ok0sauT29AekDtjgrtx2K
XdN7LDvZLpi069YejlTRYfiZjHtWJ+3Af37mAs+36FmpPl2/CRG/ynuoIq8EluTewUn0MXe42MZl
glNLNM6+RPDMfzBin+D0p9qcDjO4wfzV41Tjp+KakWZ9MKcUfE2cfVgXc4tLRFJjc45EPu9hWhpY
J6E/RnLC5wSEsSFCDxbCxBUfJPs2OFbzT1dic5AF0B6k+HJek/ZwW4M8IVkX8Jg2lSYr60U/A6oN
pWfyEILzGacf/6CJN1e6fQoc6Bb8r4oaqpKIWMUFUV/7g8fNdh/OXvy2I9dlOS8af+Ld8eTXZRNT
Y5Hv95vpgMLdZ1hDFb/As326LdZyluFfmPxYEkm/sRho2DumszlZE4zLvc4us/PAaQe8dMrfn2st
Kwx+0d0HwBWGgRXuVEHrdyLUKA+Pz7gJbOcbVQEy1a4da/8lAIutrnWah5oPaxaB5393lOISrwMC
q9GuSEwtKF/moNoZqfmVKj670tppawLApHwjFZv7HfxS1WJnY5f4E/rAa6QYQy7+z9AFXOif7APJ
p2JjyIzCsyHZdm9rbXPtQVI+WQVo8kDyD7oMT0kDbOebN09RiLi4fRAWfDPpzETmMnvS3EA/dV68
+veQQ6JH9DtMseb8mGyN1Tkr6Lgi73pkTtjEoNl+d+qpiyhhOVa94feZqZ2U+FrmVp0rT6peEnXs
ei6OBl9fhogHMnrDl0hYwCl6I+LnBxyNWknuXToS3bYORTUXzdaakjBKcsj/IaivRKYFfz7Qredl
5YjQz7F5geZPApGk5s8LUghuhJdwhIAccOkWDdAxd6ISrYEiIIoceFrmrc2A1CQTcQSLK96oT08n
1mPY59xhxfohU+XulClachb4ndWDucJqCJpaq72XQjD9E/15HY5mSFNiRcSg80IBCeBqq3VrBNU4
H4A9lLnZjXx5yPMUaXCzBSz9Wbe5b1ZF9w9rF0ZypE9ndxtsQE/T2NgipGqA0G1Lde/93hKFMFg2
SdrleJ6Y4ROPJgHmSMvS73STQg5+gkWNaaRpl7lXzSqNiYI8NgWOOTBxvK2VlKfeH/Ik/xlWoOyp
bS3gayvKLth6YsQbGHL16kSfKpIWfuAHABdmDlv+Ucqx0xAurXgk0GimTYUjmHl87w+KzPfFu6Fc
eLGn80v4NYgMdw0Ffb14VqFdl8ia9xW8k+yhDVB3qAxs6mRTbXsnnD30TiLN8i+zk/Q809g6uh2l
aBRROVWL7sB/BFLJLbBqF0CIbf+IfZcTIYJXVUEiKoUl39/OGPuaPrX87fZX94U8rCxP54edbgX8
GSKWtiNkEej6IMScEZSOupxpJ69PRkYLSHJMukCvH9NE/OKvkChfDX4g4NDRG4lJbcM43VxeFGsB
Q7B4niicFdrgOikai4EVIx1e8htQ5/9jmOB50CN3Nf1tlAqeWw7CqfPzXBsasfMZ5uEdoO3Lx9QA
6K0wIcw770qQ1pyVUq82wmgBykCUy0UJi+qQwuAX68umNZVtRIkQTye0yWq8zo5wGyIuYmIXxDl3
d1thUGcvfHYy6/6IkQyZtXk+IZu6ast5Osn9UEcARbiha19lpZ75sumJIXCioNoDpdKq2uY6AIsX
TZbRnJ9bO0xOFdIzgRjw5WmJMmd3uytlfqf0e59rgVAeLi/l1JmAxdMzb446SK+cB+nbZ50iFjVD
if1OrTbrWVK5Wml+yqYA4onSfpHBCJyHXxdsiv0z9Dei0xe2aWK0vdFwdZwVDuw0ZrMwgycKyFuK
ioDGMbcnqajs3PDPEK+XL5401lEiKAlRTBZob91uMQJVtcNurqeygu4apVk8Mq+B0a1LO9Hbmpp2
dqW10DYvDRryxM946c2Cc79mpAgw4jcHirC3NRT4q7o0CfdtSwogyb5zo+9h6P5E6TG6JLoNBXGU
945O6e2PpYJQyCe1IypdI1g1NG1kHrt3+6xXAzpz69+GRh0fTxLVSlfY8jx1i8RgWuRguuBKts/F
q/Td8/r3WmURTdISzQQGDaY1PwP09jcUn3xhLOHDFsogyswzar1LTidN4N1NdZvhFbeG+CwXAXo3
jT6yGZC06cqVJ+m/YG/0FnMKcrYnP5qE2nGVXNYQri6bwIRmiNoP86mVLDYNupvGewSJyuj5kHDh
o/1PGNJa2eBQeFpl54J8AzQfaU6Pq+fMKwODdeUaxWn6MVQHiMQTEJXZ4zXDWtSBRmKliUZqaXSn
D380Zur/XhMScLruMrUrl8KWcnKenPP9wCpRJpShslTMCJeguvgEO3aMQ6FPq7SvqQgJ4UKr/I+x
duC32cTZZdBANn36XX2iJOZ8SPpYW5+8zNjJlAINIIbQvHoRvQXobtSFv+iCZlylv07bsM0QsHwI
/g4n64VgMD5/TEOdonlR9J5w01hsuDpzn2N5jHxO2LT+cmK2FHgtnYbKoK2Iiw5MWgHChjGRvrmW
TSklebBGD1n8ENnrNi+ue0/yZE+MhApmvkOtvNaFv7z0vaPDgrY08T1mLbZKnSdfB4iYPa+KyKLV
pdRAATkGeKrSt48JcX5v9Q7q0U6AGsB8qdV/O8XCxGzq5FCyT3p/enaxbKGkqsnFUg/ybq2GBbfh
P8F1NBTIwo18Zftnln/3mp2uYdDc0jTbTPLb7ZGzm6FNLDxsZEPqPd3pfRoATC0Guvr6FGHcRXXV
9u2gzzxy+7GdB7QV6bQAxhuSVXqS1Q6167MUGOtVXlVxuM+MDjuXB8agbkhZ9CiNL1N71HKG8fMK
ryxRk+xhlRlZlS+ujHAaJurgRygRgd+FS32nKVlUY8fi7793KROcYaCkO7mpwbkhrx9dFMAqgVKf
10xAPAQa0WtdIkxxrqPayRyBszaPjUD/3kpmflqC5o4Xnh487FYBZQKZCKoKojKs5KzQ7jlNrRrP
443UHGRZILkkAJ5qJp0rGlwZas35jg5N5qIDFkgNF8tY+aXlufdEhvDlCBIGV7DtFL98T6PN345q
bOV/l5BMBX1kaijeRjjslNUk7o0uYJYMvHWFeCxliHE3xSoAStwh18bFlw6S7I8PV5BSFrgBKxGR
sGJrhiacamJhCOdQ/zf/Yglj+Eabkc8aY/zBgcUoK8kbTOvlI+Oe0zU7oBvx5T+CVtBjkj9O71j5
Eg0vb7H3bSFvJGf/unOaHsCdoLGxWT08H90M9LLtjsrEqFbkFftcKKxOAkw9bu6npMwPg++lZo/s
aWRN3+drE50pQ2DcyCBc1PAgCR0nES/8kevxZInXMBrKv1G35Jr9YkapbxV225s4jb1FUDpzUUKR
11cHaF+XilhdNXWTEU/wKJ3xdniOAjrLCinzKdJIcpIPlGhBgWZtasVxoH7ghSYnQ0Gn4gcLfX/d
PGysHdDNaGdA5i6+BuWUA422VplRf3uyE1CdAQg6Tyd8v8ETE2sk3/GhVref5zRxPFZLz3XSw918
2lJEw5O1aohk3fiWwMd3x9kGuEbKPVTanUU6RjNYrhcaB4R2ZO8uHlAPD6o8kTmOBTSEucqOelT/
xaW8utmxQoaD7LRyRa0gtxL/XAf8Y6oyjh8tQ/fxOJGTT1r5uLmlx7wh1zDBUIo9J+G/A/8wb0vy
MtZAuZJLrDJGhCswVa/nHV6E2xBJwYD0T9DGx1kJt3PcEqoEF/CTkofrZLYnUmvRJcFB4WslSCkM
+Op6alruQtRnvXQJhzfK0fTCPQx/LcWaeWozkgqx7x78XN4rC/OjdmYQxlGHPbS5Ho/GLTFIPPm+
2Kyqi8fjM/u4PACNMOUUi5WqVKGogyzIOsfN21Gtu1TcILn7qEx402RPa+1kuFXustzxg7/5NdNh
WakdGL8FLWjngZ35TAx5wLMzlOo5ESCihYDruk8AhKpDybeeraEynxISvYj5z1oNA2SvII7Thcn/
k4jy3xjvs7Y36m4sCA+H2DLRXpaF61lDUlPLtimspuvKkSEM6etCvmvUmZEd70ycLvoyU7jXUkYd
Zme8un6Kv+dQUT7eR0nmfLpf6Ob+wRAW69PHXgN6HPdN7Zc9TfVatzUZ6+oTqQ0yIZrze9tDk23E
neC+vC6uEZX/FW6u9jbv2izWnxzoXaYNnVlyeQbXpbOQwAn5fSHrcfyK9BbOxE0HNNP1EUBapubC
2H4I7uINGOFPcvwOPXD8n5p/JbBsi21as/7iAKfSx6etgn9KiiIvZXlVwvB94IEtUmVIXHv+dcxE
70amO97oqdrKF18+elwVVf2jsymlaD/bXanwOyfYPVqD9Vkqmw5fC/qXAtqhMhhms0Wj4jEfOeBy
I3R3qyhNGafM/IGH4VpI+6ZkXUEifEQ/SlXroi607DB70yPdPap+GRqNxTIUVTJHliP+tE4HBYds
YnNJOz9ujsKTM5Jw2Nin3KnUyKor0w7rviPumHq7+baWEtVK23FzjnfD5iZ9edBd+mAXeIVNV9pP
GhUhdwNaibCdlqxLqP4FTM4weI01gdU1+O0P963PVZLaRV3SJlgWDco+bhnwCdFhGmDg7JL+IGf6
qWRjjEI3/xqpJWoTJRg86f1NIN5sSPxir/JS5TigZNO1F8+jH84uFi1Z98EysCv2oeaEeqoEKdsN
NUwnaJX458rIxJHvMJvfya2vpiEWsRQorOD7zilhiyEOnq0xJU6noo5MtM4QnaHYIcNCV0YrB7DL
hEpnSvXyyPzEtW4IT2qxAjHNDZdW3Cz9mUr+T3TmvytMUvRbVo/QtfQg+IVLsADEN27vN/xN8iAH
1SD7cdAkAvXts72Yo6NhX/TUh67EXlGKFz3BsknmEePwAqEkfSMMBwsDAiqKKsjlC8STkTMx6nle
RTcczdJ2lOwiN4Y6Mk3IVnfmsUb+o9nquuWkkXXiAOXlSi1RQjX4URuFeUWixWIslip9/HAdUJVP
In6qGFBfolxOOMpsa0cHdRqaddq2BAwJ8mhD8comoax5q2TyL7sFfQ/RKRQK4eqLOY2QhJKk7Lec
i3buPmMyohsiTUqei/+uYXsQQyxrjykuMv3NnjHzOoTSo7DvDlFr/FhNXwmBHipcdEymk2Km/jJt
cCEQgrqb0at7dmqEpVQxNCSGrok5/2moPDvn8QfldYQ5ldOQYh+JqB3tKNmJ3TiDZ1kmsvL/yw+m
BbEUTbWRDtSpd2QXaxFX1909wrxIUxm3rManCi9pGsbILy2ioI+rzhP8tnZf2avQK1HlNO8AOXov
rpoWSOAU2QWtvdQpxFzqPpqKlBoYvD8lRlGRAsT8dXvAa4crV3mQkTRMXrTIWSB44KTdQ1D618Tj
hHPlyWGYpDwwFbq0FyzqMB2eTHWpAfFFNQvKQggUOcxgZYset63MsSotSeIZYPisb3yHyhtJD2by
zfAyEJeeEDcOdghFTR9E3kFG5u1t455v8FdoPL4tLX3rU74Y9XEbujTY4SuMLy9kS4U1W8TM539q
8qtkED1uDTP/Q7OMYNZSlP1Vv4+i3eSZOgDWDgV9Ii9Bbz6ZSpQ5V7GSkxLyklldituGnYKDviXc
w1GtqlpR5IdT2bLwUSguxxTA9tWRvPVQAj+lVSEaXzWD05zK7eBxc2ULqUy2CQexnuzQ2ydPrb/y
2PR0WOl564KymcnjCSp2UoAO07TQYD+g/tJ8JTzsZ/INeHTJGGmD9up+U/KEn2oPj6i9rUQ6oIqd
IXcKuNp1Qn2ks1PGMY6tZWTakeubf8TZzpN3ZBv8SGqz43LP1Iy6qtnEDMsyybdehK+UDcbqz+CT
6oGL6+wLM44bAEEojOkubREERZ7b+yfNVl2grAqbe33hyjvvs045NaKTCFt6mlR5FJWOtTdlXwet
eKszLz+UwsFZneYkY/0j8EbACBl2d2WDv8wdEnzu9ukNNeaqFdU80PJt6wRhjma5DBoczEryi2xr
7ZSPQ9ZShKnWD/gAfp5QGEaS9e21b80M/QP8Y6Bm2Fs9L2SrGaPPxgc/uEB+e/1BHvjTYI4G6EAF
FxzAc2JriYHr2zPIqOayCPChTjuI6hbvHq15XBh8sdZpSvtUVDJid1TyGNQrhvpxCjgCIBaXUm16
KRzskoZlssVoOF+1nQ689v0ZF8044EzPjLvDKxZCh+jUObuYqJbSIHGIfeBB4izc+I7QiwGE3dvT
920NV51MLfn3TGhA7MsI+pd/clm29/jLC2WVOP+CiAMPD+f3rFZEOHBErte2u5DLrOAiENmjajQF
ogeaie1S20bxqHZtTt9HWHvjK8Q1MI096kQhgi/5K9QqCJ0+jp4riZfu1XhHPuJss0ePhTrvoFfU
s5DbtPPm/aUJjAxRAdljalQdP6teAtIiO7MGG4lyde2wCO8FglmYogHbu7p3zOlVPzTxm7aUGtft
2oThYswa+dYnBbApqSO7I5Hon/LElHNaVcK4o8lU3/ljEppkbw2tMwIEdslA7zTB8afvMHVLHsbB
igP5JepYCtQ6b6j3HbJJSX+pFh5JtmWVVJiqBdS138310cNwSeL3ci/Hk+x09MlwssSa16y8iR0X
sl1W8aQLDIa6a937VJCd3r/63hzA5LIIwuTVjs76L05F9CRYwY4DBIBh10vVlvwhYgu4OyWVESRp
y76asUfPYaEYv2nGmVchkqdg4F1WTKYbHdoWd6QvX306RG+17zkmVbDqRkGZ3VsY+6CAB6q5VfWa
zqLyNHNvwTCUDUnh+lYxDbdv6xNDjl7OUOlFqLKFbg8GsvFADjSpuDs2NG9QB2ldVmeHVqicIxHx
IKTFoVB9ZuwCSTirRKRxbV/7uoHqiwer8wCRuC5Zqgfs/RX8zkzgJoy9yhTyILVLY/UUv8rip4V/
PmGjpnDJsaum6qCqAIgiMmpISukNh+ZLun+iNes3U1BSQSXDwXHIBDVfNdNe1qVWAlTseOdLWBrZ
kKhiVPWhOMx4VFT4Y8yDYzOpxc4S3jQjo5CCQMm29bpl6zuoPTeeEFna/+NXL7Wilhza+Ck+NeJS
HoU34ncrN8A/jZ1xlyjYO/KmVjKrKR3QecmAxVMJfZmyVqKXdzoFlqqeIb8ZWpv8g5Kko4Uu+b+r
n1c+9Bd+qd3b9pXoLZznFeI0Jzw1+QrCHvSsJwOMlIP60PBJFl6FexclDU2YXJAI4KAd549Sn8b6
3zlUdYJmM9n5p5ad/FuFSogvR3QQM/4uB4uSoNIV0NBZE32sVc1GooYI6ygD6CFA6Wm3vISs6Tdz
ErhUvmmY0K1JREwMqnoCD2ixaLHiM+sUwAH+/0lI0mj5YDc53b9DL3FcLUYg1yAUQn63T3piJgB7
JYuhQ3F73x+gsGje7WzTXEOPTgI9SFasBgaRgRi+6IBL3baK4tY08kMpVh4fdcdeVvNwrflf91xC
fUag6XrKa9h0j4X3ldIUN1QOHy3YcOjhxIsmNm1EtbKHihyEA2ni0VEzHYx+Ad96vAsoeOBMyOiy
FgK7jvE+z5E0G9MA1mGmX2ZK/9pRvrh7zrAyuZNiVlLUq434m4cP4Z/bCdpKWdwdFgmgwFykDl58
tD+9znN0bjKybJT0JA/ZCdwVMy+3EGaakDnMZed25i3KvHi58S3wVe38QeWQjdSEuL7XwLelhWQs
8lOI1za/Eukh14tkGkouoArGwttt65ZGNFk5hJjOm+5FOVMzCIKJGbJqb7RFFc3AjPncZ8sW0vme
s5myHb0J1cSUOEHSGx3tMEodXF39KSblFTn/Mi3ciiPiUjM+HZrW4R+PE0oRUmmsfavKP1c9hdQ5
liZdpYpDHPuKCiTai/c7fJwviDkhkw6UD2zEvU/oLjkKl0ely/VOLFOEh38ifjiYodSasUAiYYMs
1bMUpZiQthAoc0hZjSreMWXeiTlT3jEfiu+v7QakqfyIh8QeMhW3EiDrJBTGD4x9vzgHOubPumho
8ZoVnxuUNR1PxTJUYL5czX05fa68NDzVF8ErL7yLE90soIfLudlmA3zSVLuhD5t5CzrpJQVwnX4P
7Y4ArJ/UDUxD1NJUkwBxku7mTw3QXXxJXME2aoNcV58w+k3nuzP8TTiozxlFAyvS/kiOEcL48XmA
d3uzZ2SPdLChMSJbKn4PhopbmEANeNtCyp/1rWGNgU6q5vpfcEyQuqQUUahx7zXZ7AAX4YwrJjZh
vtQckvVpB29WYgr3PwJ9BMJgPAYxTzByEWnFcbk1y6sq8MNc8lrc8GRbew8zwOGQdXzG/+Zzg7Lo
44nQG2elvMhW7UMpq5HU5ZPhqXrQcuwDmxNbRcD/+ktixpjgpbZmsCHw3Yafl1iW23xBZ0lfIF2l
tU+rug4hbnGyN47HX6j3lC/H4OWykX4QIGVQQdDWYPpw2oJEGmRGOzvcgQqmnNARyMZF6UW7jHGP
LrzkSYhy2VPQFJ6edmrQqLBCPeo34KXk17B6Es2UNIQ3nh1i1vp8skb2ZFf+4fbHRgottcDKPc60
1jIsuNDXInYb1apZdSRT+of8wBX9Ud6rhaV+/XQyyWylraT5U8EyNhx3uw9dCNyzwyjr2J21woYQ
h5VyugN17QZlnNJPz1bQgvXyK8wrJyLfmrt3OHCLGgrCB90/Cl7PJ9HuFvrB4PfzHWReGg7ZTE+8
17FWjEVscrfSvBa/tROxVORadKDwA+Wg+wjMi3rmWHRNbaLjMS7tKXRIaguFWTkTtrkEJVdW2Rek
ThOg4H6UdSIPXaPy4m0UGcK4yEfZccMmnsGA9317G43U0hIFtvETE+M5EVGLFlyV0y4Y4Yz8DI+3
21WJ1yYxSs0thszN8x1vqdrMuaU1MVD8RrXxwWbtCFFW1P+amd385OhOHvinVakHxgc4Tda8p09U
yF3WiuVU8zM+Mono2LUK+nX6phOsRXOlCerCh+AhPFWk6NqOvqgJGKJ6drtbExUXf+HKkshr/tW9
ZHWi11WX0JHLPfaVpocmrxwl1RZy8stw3Y3DCaVbuT79yYD0wHHxxzylgTs1Ma47CdIzDVftXAvw
xQVOKRZUoxFsISC47Gr563zEO4MigJufnMFLfYSghFFEDtUE57mdf4RhkTT4c5m+Ft6FQ1Tq/dPv
7gl5GsK+s3ub2H4czjbeyWGmwjc7YcOYn4BDUk/J+iZ2b534yzWhiGxv6UoWCP1M8Utuf6YTqDBZ
N4Xw69ZSIIIjAb6iRzmwehYlJJDURu1ubW0UOnJcrYjRHrKhZajkK6FkbHBTYLRNjdjd797qDaDF
+MHBbLjKz7SkYuiI0KfUltvE1ZbXfKPZrfMDPD2/FshXJi0FCT0BjZ8O+FWBWYFMaMAfM6l2Dd7Y
6zJjHjukQ0YmlWTQRLlljeV4w1PXJjy4eCWVoe1CZHXX1i3aPbMctS1aJ5TprOYT9HreRSTMEsy0
HyGFjFIs6dhSnycUM+VKpCI3wzlDIp0MWO4GheWhKqZCYXy5ILKNQyCMDacve3vF2O86aV/I3IL9
xxLSeHTey/gd9kaBa8E9631TtVlK2+co7noyfz/HgoLSgLhxR694GjG4+rKNeuCstoKrCQtF/fEe
YlqYOXPYjEpsiaWHF7aAeBWF6rq/oDLt6X9oLqD2Sw3GDOXsgTvx/eplCEVCmU9pfOQrutrYuDyZ
AlpqDCWJByiqnleIW7yVTLiMWkuCs9FXLIQ72PJwMe1pASj964gPrFfuxrIbRkvBEioOG99Ko/Kj
8oOM0yx/vIFDhDb014rQWoIpJ0YzR6gQFaKeA9AB7miTVdzdaFFck/RjBxHqs9cBUK4ARfCsRxp3
t0utIl3WNV1kMMgLMQYbx0wxglDg8lmNd3winc6XcdIdhC0dgz/a7ZE2Jy8W9sMHosaLL3Ju3Cod
DGwE0v2j5Wm8LVvpWD3wxIKUul+G2mhEvwWlD3vNWQuht2JoTp+itOSHHHgYziIgTyFDfz4V9A4o
U23JYFHpGznz/jTdD0otPSbhzxby63P0N15vTmzL4rKcZpFQzLfTnDik5ZS+BvQaw4ukQ86ste/F
0L/24wiUilVeQ6eDv3V8uiiio6Q7ELczYwqSQIYGwCNiFvaVm0tyafTRnFQlAxRcHAenJmm69W/i
CQDU2eWrhzBfrVx730Uy/4mAu/47XsiacyMHrISnaisQcO+KwP866NxDCsO5l9UvwsjEpkIj+ZtV
R+tTrvVMkcFNj0HIZGS0DfvoXgLYM4wIELp3HlIkXx9/FtYm+0oi34c0pXRM0+ZAKB7DbqdNfnJO
W9K84EcEMEzRTGHMFQW9LmiPGJ0fd8+DPcyugNoz5GlB8mrxFfpQF4FEOA/TVuBUVrRilTMkWi2K
YT19I2ERprK6LdBuyUDChyhZBSZdGzg+ZLdgvK6KQHMMdt09vNuQl+QpNqlgzYcdpyIm3VfE0fUX
53/xBavm2tcNZpPkmBXjZauPesJip6dzvwXsKEo4pRghA1iJbN9vtSQKpLhqCrVAQU52Yzw/mUA3
6MVm024aTHws//uxHih7ZI+d56gV7ujKunr0LFpynljQQfFBMIwFPY3bgmqMbi1AY2wYyytWLJTs
bUIsk8R1bXf5vimpHn95sdotodTbtKBju1k1FgS5FESDH+d1ObAioob2WLgT34GVMotCx9a9mYqc
ZYrstGJpVUPlhM1NMCksBYICPRXNJiq3f1yo89yc8Q15pbXfyAnxcZFk7Yg0hjI+vBQ+czgaQ5aP
Ifo8Ia/xg6oz4R8IZC+WQjNqH8asZkNFQ/7zJVPD0v4yw0xrX86+aqpL9y6I08qobAAitEU8AVeh
8iPY16cQCHUSCWPK4BW3HQbKIKtxZH5NI+NpqckksgyMwlo/22ulb36Mm5u45h6ZlIzFPq0dSMtx
woN8zqXuGOukfWWABQuTe5D5UZowE8i9Ctc3RR53kBsBRvqj/Mnf48SsSP9FE6y1ZYMU0Wk9tXp2
SAkB7FmEbuAM/NPkf6l2LqiNf3H2B0BUpbVL8oendEcRQ8WpP1UuHlWy9wSWg9efm+YzhJZAzoCV
EgbUssxHHeuuTAzB08IWQVnRGmTwOtmjtppObC/BfKnu67mQ3UwLCULYxO1graUIAvrUNaDRWCUJ
/kOWQS/pZVO58BO9UE/1jgvxVz5d8W/QWO9wIRSJIFFauihac4s4BJeIC3qNySw7rUiwPvpyfGwf
TDAoVIZ4+Su9/erJ7m9JOSx8pQaAKLPkQWWMlDPXy7Ryjd70W+UAT6zk9eZbAfnauaWtF7pP4+hF
Q8UA7R+PP70mH57kgYljnQyXMvtnJ++RXMC+GmY6rGjCNcxmwpYMIUE7DsrtxVCjm8/65AZqoJUn
GIfgsUpor8KxmJqHgZRJN9XPsLSNNREIBRIjbSXCJribEuT5AfKHxMsymuhlaL6wyxWNgkbRitSn
eaD51JG9TqUlwRD//aGB+yPUs+K6CrMdTw6QQHum7I34k5q061lq81VvVJC5lNzMDZnDHVvdxZls
zId1F16YWeWp0oIM0rAdJ9F/wlmpwD5qDyjY9gdk6y4clIkqrXJ5EN2K8IJ+KNPReE1QolGmUlfN
pCSKX3N/iFeQ1Js9f0TVJn3BZa8uArVdffJTT1Vxss8YyC/YCb/EF9kuUd8Mj2BgD+iD3nts4a5r
r5PqyLnNkKSnp5QiJhSnWGRk6K+F4Fe1bEjBLPefJDqV2Zo6FsXRN7RNBpUCtInqRhMqD6fA9ceo
T7OZXu51tkHlSOWLOnyT3EJXRYX9rsbmtoG/RFnnXJZT7vPP5yfuaHzrbzodvkdHNSSRJ2reoM91
jRGag3yWXH2avLh0Z3JRO3Px23HW54BnucodL8GaJ0x7hrd23YsSRjEugmPSzjZhO4OXRO5/KtuT
ANhys50+84/J5cWOJHiXXFSKJfbexM/IwFud7LdljkCvPVdd2TmMTfVwJ7L3k6KPLWAXiw3tunjA
HUhJlBq90zgc1TC/f1YSStYYCYWiBy1MTEFrlZGKdDpesUJVFlyXzfhh1It07aeWhdTNfaxDB96P
ifWZ6snB3qoTl2RVW8mt0HQFT0MAtEaKfLjhQGEGoO8u8U5QugKTah0IL7S+15Ep7Vbgm6VBvu6G
p/2TC1etf06KkXvGUAxqakCHLAzdKMxrdQu9S8gWNlGh+t4WbXq9mOsna+pHEXyjmH28sBS9RAU+
ExSTEYXvySEhVTOH05Agn5rUK2GWpgdHdGR7cGD4F2b20r8UkxifXzw1V2l7R0VhQ8msZd13Oc3d
twNVwzsYa2y9ddObKzRcgEH2I+VCYx7cwKM3EcCOvIcPUdsHDZQuI7BtDqpToInzumytT8NskcUZ
eXEYEC54RN7tmjL8kENjThJ878sNy+Sk+U/P8FG97YtXihODOS8HmKpsnaIOgjVBmSCRceqk55lC
Wqg+i7m63pg7p1UPLh9D3jn0RoqSURlaopk/7DsR89BhD++MWsfHFhGn+mJ2OxhYiKZ/dL+xuPCK
/S41gFRE510tgH9Q+yIa3FDBBmUUa/62mxC1tFTLBRctL0jKsXkzzPU75U5uv+tZr4681rttD0l7
TrVpK0i2KBofzjJPgbR+WkY5Ppg8WXU4ICnaewdAdygmwZkDdExrmsuu71TTV7V5t2qc8AB+Llq2
c5KePQPpJPafZFmGtB9rWyEe9ctUa6VlQGkDLza1d6bTTbqq74Ty/MFESMI/ADxIqqMNypI4QkJQ
iU+burPLA+dsVN8BmxUBZZalFrkYVgBSdu5pyhcwcW7Et8/DHk9RTbzEFCH5+rFQEG6pBJrDlGwr
G2VcuNA30HKXnLgZEvZVqYCp6hHdYgcjLW967KZX0CMn3mMD6yupyzVIqKEGVNeXQHV5w5ifQiwY
p5igivAeQDq7v8OQTu/QAf1FUNfHcBJJ/xTiTOCJ6BEXcY/UfqacMaHCQEBaqQ8gSnL6uxnu4/Kb
jMZM7lxsM4IRyhvOqSVJRCZUASZryhelPVqx7kXV9KOtC94ivuyHYQNpn1T7srxDVPhFk999r9D7
i7eZy42YPZhh3ItTtDNBH08Ena8W4p0KmG3dWxZD5T/gUbUla0knY/39+7V5ZxXkWt+CaGJBYrMo
j8HjfrV2qanaaZrFU+POt6SqzjQULUl8Fc6udURvSCjhUZ3FuE/4A0Kdkmoy/Hx/luvKzcLtbYr0
xhNQorSyuPVlovsnpdayCnPsdsim8CnhGqCphdvjHe6LcFpAH+fajcTBtqK28NZmkOQXdEqx5gsv
BjF/tcS9hSOvhZhdx1pfUWktPetSzViALygS6VB1sM+zPgg3aWcJ1GRv9IZ7OQods7T44JvOHNmh
eHJEMWF0Sj4Ibs37HX/Rn/YaJscSZ+If+/FzvNpzgXDjiI+DKMQdc3wiVgb7UWZGrUz8AIiB4atV
gJVc6Tcj1v3xRkmUYEE5CB8Ko887KtIPP4bJW+0wt3PHCgWCIY7u8nesvbbL7cX3UGlUnDcsAo+M
EUrBFnYPoH8X3gM1db6eftt6dWiNRM1MBACl316yQmGBiQQC3jWVAUfYVxojJ6BTh4J8626aqFIk
bHWYeGykxpnNPEJKcmptVkero+ht+TkrPKsFdcQ/z2atlsU02BdSCeNNjXfM2WaH5CIfJTU3SGBq
q2MsKY/nHtSYGsxv8h7YMEjS59kOATILJ4oULj0+3do7rqNxAKXR9eFhmEiMW3Y/xOARqkSZYghU
ZkQ+tOcmQBd8fmzes+PFGU8XRZvRjIW118uieIsvUd8T9k6mFAIns6v934mZMEHA2uRtOxibxdHZ
DRr1fhZcUW5KwD3In4U4Ppy0pFSx5gej6pWHta0p22s1KoYVIxfrN+BfnnRZg5rUU7Rm/+Xv99i6
mH6YDCzO0bYsQhSRb+/Kocx8z19MX2FV9iGIHkZmzIicdx7O+Fjq7iWyvisZ7aHLPcWex9908pI4
2nxdkSe+iCprjzhDfaycbmdFp2k2dG3K+l4Wf6thYa4QMVRscj70XzUCY5muc8nmcwtkFaYldEuE
Et8KEgaBbJikZWH/EUFYMqb5FF+jcmvPDLF0K5uF0l0F7Fs1D11uThtwQfeU8fzP0pZIaOTWjvhI
O1dhlc8KAC/xOSq+ZNaeVbnF4xpTeysBfhQyYjEaZKdIC4z0guRUO0/HrTLEbR9+hRXmnYkJOFCX
6b1AsRkcXEGBZI1HbZQK5KaLXj4p5uefvwCHRFp9K2nhCg4/cC8f0CdUu/NZU3EGnhnPOtAZvG8/
/Mk8LSnRCxz6cFYAEw0EmgwW3qtPeqIGRdEdJXZ/Vh2NHusATcZxN29A6ngKDKLafYb2NqRPv6Fj
q0q0DOWS2uxsyIUAvzxJSigttPrvP/TQoAdsbp6wq5iYtQA40ompeHGa8jF0RHiO/B8DLx4lcR4O
nn5gcUB8Bm5RkinWbQ+EAuRAxKiBgPk641aT80Z2pqWVLrEa3r+D6P5sazyp2IjFhvMEpxdKkSgr
h6Rx7ru16seok2fCJqDW+BAKN3m8rBAO7Bkvs3yi9sxpPFFi8A1FQYInrvyG7sUi/53w4J+t8dxy
U4GWox7wQRxviNjvvuNz4nEHTkwhRva+1Zaigu/2ejCVCrjihZmGmJpVPDEQwsZRPQsIFNyuF5Sz
IrXJUZxDBcD4R9xK8IibhoyQV8xwuHs3ud8GgUwGvU240d0+QD5+O0cuRBw1VGwN2XKWw7qFYP3u
HVDe8Bj3HBDxRCwZmbgpkpycBayn2Wp3OG12g72gXyeWuaFwo9axjPCNXKtXJzc+D/BGeEYvPnV2
dBEuRwgu/DGYf8yJaf63aClDVO95fkff6OuNJ++bVh2y64U7sEotw6zK3byVX4hMdjjqrBwq8nKW
xJ2iGvkIpuMEeE18NjQNgVMzrIhNBT6VV7ZTxjFsyHW7/a+So6EiurJKThkHd6pf5ZZkft4N7MJ/
CLeUYetJSODesMwTaJWerKBceEgCiC0lH++ft8vGvLWsmJsw7GSBFONJn9avBqDJtiZYS7yhOolu
votnl6tLPkd6ZlDid0L/hdib5Tbt5GpG8LTM0ich1WzUT9DzZir1KiOAyMhrOwxStztkCYnIBSJH
xJNfORGmgTP+PVKwhYFRNwuoknhxVZcD5xO3pgEuuekSTk5mlElseS9ZUBQWZ7yhPU9ONywcBC6n
KEKzRLXYDcjMxEipwFltCEMOIfCtlviNwoLkajhgxQGbxPkY/EW1SSrb4UfAuXvjcx6q3/Tuv/28
uQMA4lt6QNDPVp982TO+IMr/bQS5Y8uzWUt8ajohrXLFhKCYWhE4oSMPqvRsrMDVi6uu9woSonn0
S7QgyuZRXXfmmzfSoD1p1uwA13LGL1nKxWikXFVMkcSHtMU4m0Mu91QR9jJQInx787zs48elya84
MVUX/HEGpQdTrbmR6bHXcaUvAwRa0+bswvFb7Yvmae/c0MrNgElRQ8IIOXzSdcemaDzk9JUqBSiu
cIYifRv1hO7k7cWNnwpDcOTJFPnmlL5zLpG4AGM4QhsksJrGkhFDNuxIrbx6C9/i2NwOD59V5Fr4
YlEmwgFX/z4MZpHH51nkfz9LkqHSGGenVEcPgNpkdTIgyzwfECV2vLSKoz1DIkQ/zoK4FuTzwE05
BRyhDNfO26oheVvKnCgtd2pl184mF2fG5i7X5eKZ3qK+jaksHFQAsd+1PUw8Ye8YKUAu9tsmGZYr
phr7fqGt0H/KQR0hAUtJWl1/vOlHFhHtZf3yesKVvfUXfTIihXGFJzmW7RK6NIzAd1/uumZjbTrO
SISvSDIOfu9+B47Sn3UtCfL1jrhGtACaIHJJW3tV+5kLeKP0yd2mpjyrqQM+HSlaze8jUOs0/9FU
1rFcXABYhu51SKHam8bsCxQh0WPrUC8bughcIMUKu0TubVVDUTh/xeQLK0YGYB0VgOURfF9yqETW
782tpJ5pqhARyx8cpw9Gyjw4XBOODdrLmjdu2KQKlkf7TcAjy9Gvx7scZKzImxS0z7YZm0jkrMsM
HsD4Q710ESd3gza7ndEF4MLUHvSiqWCB8LqsFgrgXvgTPlXJGt6TSJEFjkfjg8HZwoENcBrJrvze
vofDhZAUdwW+XwauQa1ypuo/C2JMZVnzTUHmJmb8ahb1SqM/253EKkjNGhw8o+Gyllx0SIfo33qj
3noZ4+eeYERMBP1feyJZ0bOBjsWv5HqY0EFMFFtAGVSuo2xjJyuFX8e04O9ezufouP3eZE1NwOdj
F+/FVrEYpZfpUAI2Bi/D7wJIPZgBRtOxLcQKyLj5ns8By8/Fw8jZvxVQGaLIN9HDIoeZCl5TsCsB
kiy2XMOsvUKtTd5FYn4gJU69sII3t5cyCd8mowBpkcstJhEN8kyxDyouTwzvVODJMgGMhutO7zQV
ex0kAaFj1kVpbqeYoma0vR9mar9p3Lsb1rgmyaeSKyPi+Il3HrSb5BMO7WDwvIz9HbCmjHCQ5MQ3
NqQUnRtd3gg7cfoZegJVbg7uErOHvAcamCrvUkAcOGIAwYKir0pRfMbZGTUDWN5TTutdKDnsr6rr
WjCXAGg+NtfYeK232xeYUvsiP7mv2DvicJ0kavzOzmkwzys62L+ganWeW4rmiFz8yDQu1UTGbcrT
rfJ1XnTFhfx26Ql0qqw46/9qIv9oW9mNgtJ94VbEOUpzT+IY5bx2wD9Mcu2/cPS7y8jaTES8WU1K
CbgAtNZuA/5v7ElfrXSCBDfuMClt8+ojIHKJF0vkL3O5lgqWIlRQevlPIV6/m8I3K3Y3a92jUe9u
Y4gJLjRx6gdtgrdhho+dVQPQ9A1NXIKBDsk/l5aslQ+IjVwyj8oxkM2OgAPoXSLigjy2A5vnSQXr
oGNUOxgpPFb+kTmrKiZnX/I+VVmgwM/APxkQxwHeYquH/20KlRVDaqVKL8GqQaJ0NMdeeTnt4Tya
q1mZB5cjCHh39I2z6Ayxz+lOp1bI2sXRFxzlJjsxzVaRnRVJLr8bzb5vsSCJCr6kTjuJ/RvIt2vO
6O2oAlHANxwATyKtt1ki469/kdI1KMzU4teb7OQv/TBv/3A2yy4G8TRx4NoNQE3C/K6IaSIkB7Vb
gf/lKxg4I1LYvKNNG9ThVYU/iyVcCt0l0T2/CfsjCEQJB911sWxAwNu38mOEfAhL4ft3OUEnQLPO
NnjIlqGwq2KvYAJSGzjkgcZm3RAEaKuD9yQGEEZmpvCyp5sTXkEIryBB161/r9MxOiEcg32P8205
5EF5NGI81iehYFFO33s23btJdRQoYyFEOywxRqr9B6WUhr2g4ZRCEQ2sO7g/VDIhUXithUya2W/z
55abjG1DHfIFJuyTcsuk2l6YOmGv0RIQiteycxxZ2KMpitTEY7f6NOHmQGH3qbHrK3VUDNCctzfc
N2WKSdWsZajLbQIRcjAj/LKHZndHTAEdHoryJ9sgvxa1J8rx4jvL8BlV/rQKd1PBDKn3H9ybTu2G
uhGBPNw6q9pfjekKwPhwdZHfhBDUH20K+xT8H8l+UzUrAQuHRFGCAYz+5ZxbFW5F1AonjLDQKCU8
NFhQaCTRoZuYxP2jQFg+oenr2ZCt94eVqUGiQ/9s5cidN6ysWTRw6iRbK3CbNVKX8s3wRnaw2qXI
Bz4bSSxnT0I3E3NcCXXZLg4ydC+IKEpA8rVFSu4JPIC2BRStRBiz7i/GSyrc0lnVabnk6LXTYNzG
UdmmjMam2AD7krkngKiiQXyc8DNipotOJJpS1E55O6ranT27RVFVkJtLg4DC3p91d8O1HomQwDd5
t8H4GyT8F9g0M+nFX1UQRYut9JP4Eh+qIikLTaj2S/UHQHn2gESoL3gAEjnXu4ZL9eV6/3jlXyt7
lGNS4nInE8XSRd1K3TUF4p+YS1nZIAwnK4mFyhU7T+TEKBZ3thtm+0ZR3wZvStmoYn95SY6Izg41
lSG/47Ll5x5o4x6DHfVaQIr4irU1/11dJo1OA5HAWZFwPWjbp4qo0Nb43Rr0QPEf5faHMCArqlHj
pBS0nzIsMUUPVIf+vnUtD3q2gy2/b9p4Pnw1RmWKwwv8VJqaxqNGi/m4h7z7WvHdHCCftqLXbP71
luGo1gS2AEforSTrNWSm++uoBvdKmkrh2or+gx/UDEP9DVvWGdWWslDimNQ/LwxvSC4o7KZXhaAT
CPlqMJkdIcjZfvjms4w73J0BzDjnCcPdYwcti6cez89C4Nks4abkGHwR3RqQ0Z6o46yVxLlkza+c
4AhyJeIiHv3GlnR72DGCxvY0MNiJNx4k73591mPZwLIWSqdjWXxX+MN+JBXAdGMMvJnL1g+UJ6i4
xMyrR2zwi09fefpZf03mOAFLG8yT+2Aoi/q0uB+zfwamYMtdpInOFBglWi0XO70gq2vUg2I/DycC
J596XdumV/AN8yy+pQznjrNi2dBEtnH0eA0FMv7ZKTibl/8yWk2+xhlVWkKgNmvt8cYjZfIVajS7
IoRsXqVc4tM9yqrNKt3M6XGuo9KdHBVWZOp/5/+SgST3zwDDouNw6bm73rDm0C8XtINKs6Jyd5O9
cR8MATDz8xSZsmO2PYFKr5beoXPUlriv/TJL88E8ZQFVsp4mlVX0yN/S53aXgpvDalrAxXzi6h52
v971wn5c6vwyFwrmewZ4Fg+9fg0SyzbjBijcHFejdF8KG+9x2zxDy/oneQOaKqtoMZYzKkxW1kZH
ReUe1wBB9gIwyvTDfqSeQGdVVRAJoXaSpGC09UJODKsAVKfEh2wECxW54M263bJCTta+N5JZXrHy
2/LgT1vLE2RnIwBkIdys7WH5Tbb6wPXc8wyDqStGStB63SQZ/TNgHkCftFmY6tzB7+S/v5u9U4iB
Ias4EMIlh2Q5+p03OPjkk4MOM8BoLCO4jItiNG373poBybjkUk+tcBo8krE7MOo4GzzBuRZjB03X
FdGrS1dN0KVrsi9WuPE9MTTgpqhBMJEftJ8riEHBYP3FFaCNQO7WZ4X4uaU2nUGj97Z+okud4Gne
+Pse1X69xpXvuctAVtRlgIM8GRg7ABABFhsQLj6vUiDESNUMOdrJ9r3Ev48XvFqJ6dNp3n4J+qSv
nMGux5rtnB0renX5l3W100GrkIJIDPfY1fDt6T6YQHOKSkVWaOWyoYMfDJQL5OvNkBMzUUUiRNXp
uVQY54uGSxKv3CXtCWcLoZE1+upwCfD07yODJydvKGQNxonViiMJ9IO8hbyb8+OF1TDKKjjs7dTm
4KZ4QnHGglmjzr6UxIWXseDZmBqlXDCdO06L1EdbCwDKZ2KAqZQHjIzOzy2Kr2/MHb0WGVEcfIDL
XNuf3GD8DCuALeXl0xo319Cdrzgcd6xwgGzk3n4x7X08egnL7J+UZLclEjLK1huxI+867pRLKlY4
jpY7uGPi/gGi8IczviB8dgUpJVOGoBFVEBTnofq0OBlTKAsDNHK+eT+KtrIP1vMH/Ur2dxZAWvUp
8+qGChrlqgMKanbvKWVZxty287I+gGckOfYTBB2jZGmWHu/XT2pkM2+h95a+hPY1mPiXIiTMBFNz
qe01zfAqjWcfanhb5M/+XWT/NI/F3Kr6uP0Vea9Hyq3KAKLU6ydmb73qWNj8g7heVuYVpvlIPJi5
1ZY1CHEbbRhKBjGekMDspDkwHFFb5fJFqefV3ZxtC/F9V/x8yC+F4i+gQMKXdT2KcMqYJpBAPpik
0XETPNDb/59FbltJou3H/Hr/m/ROHTdPejgMZEoWmrUOfc9J6zlgH403FKAFEkQXzca/f384uKc9
Wt6IqAE+93U8pqzXfikGJcBOQnwcGDoySDPzpNdAEitlDcK5/Pz6JHoUeiDaDUQz9ZXp6vDbt9Bk
+/SqE5nrJoC64rE+j4bus7DS5d/AXEqlj5w3ejGrRKKHrjJePn9zTl190Z7/2KuaY4yZX9pcfJPn
RIAXlK0UG84PeuM6bZkCVQ2U7n+e+c5UWhghyfq3mZo8qz4piivJMVZKpo29ciR2ZT8678XpgfBY
zToXN/wEm0sUURz1AkzipM4HXb/miuvXONSkhAk4rCI9fhkJFc8o7w8vQFNn7xRb3u4jwvENEMcZ
05XJFnwPI2tlxatL0K5NxcI8udTxsFcX7vBmLXAjVRrKNGT5gkQR2CKt4kDYZBORIsUwxA1lIQJ+
ONXBxCMtjf+UJm1qwwlDsLD3ZzXGC/LrS2ZBYnVTJURwT59FmYB5twnFMqrnY4PR80HFGWJK+U0I
VJgZjqoc1z2O9DvlW6HdshO0e52c7YNcCU69ugkjcBI4cidi8UeKPSPeaiLZOMvcRQ++u3sNFyW+
/yASiZUdMStv3UTlgmaeMQ5AZavrFl9VF0MhnGklAEa/oeTg2EYthst2e/xjlZ89nlUe9SjNiO96
FAG/yPtv3XypmNk4QWjzc0GwqdlxJ6WzYJyiSAwM1Q8H0lZ0abfg1z23wTeOESDTQlPZyKlQikv6
ryBVAmF+mCG1t6/3ReoDfvRdx+BpzySbmLAJoGsXIaTLIKfQkAEaGGyWCWr0eNuswVa6iRoYq8MD
Hurd/zM7O/gWxEQvZmUCm7hJpf4asd3qHNfvH+HatUv3JQEkNG4W8b1H+MAQorRFP4w+ACHO72hw
QkHs4QsYiMCrsxAWHaZUjzAr6ZNWij6lkHSlDnzYYd+MctU4PZY6f6XkvMDBDAAopbT/agHzXAce
qYpTSVhfQb5rwZ/yXCozDVSl0fnQ0VX0+AnIWywH/gcpfgGIh5TlNW3Ifb0lX6XSpb0+pdPeZUoy
h/1GcLAeS8s0TPNA6emEx/KwXAillCp8skP2xnYIpfq76qiSWpe5fdvJzA2eke59Fo4t3hVLKSml
9p+Mt26p2gmMYdnaHNq6W3TpI/k6QdMonKEjgk2onXlvMmu2eVvV6Tc/SGdKuhSUMx7t+nRAW6aG
H6zE6/tcBLOsUBAiAZ3lazOJjP0rbjKrbRCQ9vN4rDYU/gou6RB7h+q30VAQvtGHlj0YFgo/8sQI
b16EaVswWbnzrr/WMkHwwdV6MSZzb5Heil9GuOAAN8Rd6SVCq3uGBhTFv2aVC6COSHSJGaXNqeuf
+auTxfk0VLbaofDT7CBaDHf/2BHC0QAuUscNobUOYy99aGABZ2wH05l39QVTyoIGnMh5UxWDscZF
7oGQLiGGUCqLtsXQm/ujAbNjDIaIcSDMVbrKNbmu6V/VjHWaHir5F/Qt6HlXkE2KHdQNkunutm/G
yD195s7sMDiZVaUNWtAakSqlVkq+zkyKLPKCSGpruNYhidcvovjC/2vO4oV1EletpDzLjaF9i2R3
+/S0YjtnSYJcKtngRgC40tK7XPZndDWV5yf1aFN+ogjKVFH8pNbKNroI+CbPtxHgY6lTcXeamKCW
KmlRIwYUyHUzQZ6YAMREjTbqDimCaNBJmTxH3ux5gz9MhkvZ5ZkoVXvKsuGWPRVHEUrKRU/NUY/M
vsWZUZBBGBN5H1x+xlFgPU12JkI/1ZX2dWwPSO/7ycK8UH7GjuMQVRfEeKNVeisQFKC/EjMZA+Ds
+H3kjWUwb3gexplRhly85tZ0u4NlYd2wCnOXN4/rpSWQgpfDlr6LniTf7dsoIcRn8HSI/KYdRYIb
TTkdGHTtodjeB7q4ikk8OEv/i9iCKzgpWsSj8MaQbB0XYdmmg2B+dquNEhv30K9j8KQ+Rjp//dDO
4zRzt8tajcsNeKiHJzCIg8JZ3gGDWRl0AlF6inN8gSUVUrU+/4wxt/jOd2V/PGoeG3yohIfAB8jp
Q1Dfdtkz+84mGNxwWGvKkFZkT2MWmo9hJ94LpCfnkiiGeZCBIdQ+ewN5VsN57+h4ojS9pE2847TG
kSU5O/s2fQejnO3EZTtdp/heZUuWG43Zd6hwRlFeFBD0/AeU1BZX8EI6ovMeZewQNmNCeKbII+gD
zOMcz9epxyI3EoM1yIrmNAysbiOClQprloFn+nM4wa4rhvTAE5wP+h/21hSfsOqkbaVZyd/8KONJ
qHawqjS9QCi5XfTXqHgBMwXJww9ayD6yLtdyBF0/Pe4Y4n5bigkocCQYQ52Dy1ohCZx0j1iNV7EC
s0cPVq/6a/6A2DDb2wkHl1VV6jz9HFTsKN8yUb2c4Edo5rEqGaqMCr2gw4QUjeDugOAwfn5FjhPf
4ghjg1u7lE5LwGpEDjk7zDCbOpaUUGLuqvpEisyVkUOcLdEcRvg4ByLecUW8XQjSU0DHCqYyEQSb
fvZbOkq+sSoy6BR5rIuoLvNSuqHQUww24u/D+JegJe5v1Boj5VnF2pVfUbVH2tW2Aa0IaXSbyRL9
NMjXPnICtjL3AM+xLfo7jidje4kwNhYMWszMkYNMLuBZDbGGTUSZKiBhQ81GrZnaHDkT3CGk+rl8
HuFBSpreUkulJvYGTUnRxll5+txLrgG9h8OQmQot4Q/hQF5LKxpSUp+TGHmojgjBg0Bwo0S4ixT1
5v0cL1ANyCtqsVDRN4uEd1QZawJjqW6U3IJJEddeMCSLzRWwxqbFAi1r6pm+B+WRLurbXoslaZ1C
Q10gdxZj0ewqdXCeNNXrZSoFIeGvNyTYIK1zee9NNfsF+l5l/SkcsaFEVHVpPtyuRrtvcsLj0AG+
5evo7xjFEaimrVp6ODlRd0dDJRLP3VknKDc53nkmWnY+tlRXxLqDvVFQvr2bfYuHgSBJf/lZrN9T
nwrAvT9PBqTixg+fvP7eESs8qAAI0yXNUwiU1KHyu4Id2/9Ph5y/fLTkII5Dr4QEPm6uepPaDjPz
mZZGx7KekneO5mK9BtsfCsBONCVEbyS7i/9eS9tg1hNyqZ1L3rf3mn6BDuNuAVfyqOLY44cnPFNG
5VIpX12iGHVd5gsZR7JB9/3QuqKYVDSqznmxgO8oAkiKg7KRgd2hSzpcUAOoHy8WQnJFMw/kcND/
L5yx1tm5vsYWaagfSLdnrPCIIuWKhiR5B0D2Na/Z2C+dxyirY4qFDw+B2W1LOgx7Fyx43LgMOVo/
FBXB2+byLZovuM8X0cXg6N7DvHW1InFzW0bhVtUPef7jlTa9TGjutsDJ+Kr40IDk7BfINneGrgFT
OJJp706lJEibhi8m7C/MjW36WAYazgFHrG0DqpjZwd4K7mxyWqeMc2EEvHS2EtPFLsBQZALNNo7F
iRGAF/vHyp0tWTKeeLoB80YSygqCiPtYWeJaWufXyYGkyL63rY1NQa1LFUTKjjP2WOctzs8J6Quo
r5ZrVrxTOcXqkaTP5nAMuA5gGrS4qOTxpZKfMG3QF2OiYhJYBqewLxyJ5SEJqJuqMWixa7usEzbP
Sk1bTzQg/75a3P/jPQaqX9lsfKNz49GiG0Y/2uyD6qusbBDlxJ2d0VbgH4zNpkAfvsIaY23+G6D8
0Lq5O3YEx46z+sm40yNUl3MHOeeUOgqml/evmwR3563LHtey/egPYNp04+Nk/3FcXmWL/Cf7b0oe
z703wFrwD+6tny8ojb3Gg5H9IjjJCx3gQB443vdBqO/DhqIWM7DcOs6LOjJ/QsnMiY3uQxiY+eFS
+VmxA52jRCjlcy6hocagjsUsTp6bKB20PTMontPhE82pJ1vMvSjJcU5hTMevwAVqg6kH2NcEn0Gf
NpHVqcRl1UR4HVymE7zOdkJgOaPWUk813vBhbCLD38fxq5J90ytMkJL4hF9UAhqGpyo7cRcHeZBz
Xthprl3IazImN8RROR+yhab1R4kUfAbzVBi2dz9SrP61915cY47XVXGJ9baUU0RdnRE/83406qtX
toF5xTWuOHXXuEjGrkyNXt5Ka74YwG1Y9IKp/aP+Y0NLK9SRpBaET1+cBG/s3CJFBrk9n0Pd6cqV
VAiAx21f8yzthXqod5g6PXa6ShD62kg6Ym3nhZQ5AjJZTXQd/r0nYK1tHRJMoskghShQ+BZoDqu+
K76/LgMIWxLyHKgqWcOk5tHRFWWJSng2A96RN36/mzONgZauuP3GRMxtcdNDT9/xavftx8inGJdx
4AuGiRW6GBavWFeuQe7CRzg72sAvWxwTxIHvWKEgJqO9I4Qj6amOgBp3psbQQ4qbitn2lWDaC4Kv
ZXs93u6/KTRwIMWdOZmoDR2OMT+RUwrwPjjpGiCS1B9UfQXOHFMIPckAi2fruSMMIkDlnUruHBkM
gidL+dzjwGLux5q2/TYETfZFlayDxz8cpElRWawk1PfPp28jFBVwa3n9GxV7Rd1BcqDBaWciEufx
KekLQKOBQ1pwT4FOIbjWfWWFWd6xQTp8zTwBkjzVq9jEKfeNhfp9L7OTUE2LXfjrDRjKW2hjBYtf
lJyWxNZuB2cDrBFSYcLiyc9ThURPmXGU635klZQmcFRNATV0HKTilKK5QstiT7rWypWmyRKPji0l
maFIT6hMRFXxD3KYolm5eyvu6A2m3eTZSXbl2su9R6gfLyXbN0+RAU83WjG+If5VMe+r0ukL0Al+
ECJvvzxUWg6z7UeA0UwGC4vihYpplTAigIC+1+yQzOIsooOBI/w9bFXwIKvfjbDpCGE/6VnW/1Qj
cKkGSVkQjS/D9hd4co6wQrreKJcGzmBXax3gPn8J0CzqHTb5oBzNxK0cGPn88jt7qpI6W3mnfgS2
XUr9+K9kYSqIHd/O+BNRJ8G/P9W73+mfqJVOQaNWe1FOpdThzYw/TizUOPDEfaXEwcBKsr5zujWb
EcoUIICdCzf9Qh5cXDXVW2Dwr1T4TsEuQaw3EfIgL6LCBzLCo6pU1+pU9LKePZGa/iwPPDJKvo1e
yifY4m/hPBjYA+GeWaUb2FVqCNAkNM7aWK3AZEmpTD2uqLXVekQndAhOwEe8c9RNyQMJFuaVNLtb
AreRjZcZZIKiUmXUyYP2E8VTOshpL5I9zFMGzty59uqviIVGBSS389iLJ/f3Kix+uI0B4dHFLRKU
Ii0X6snh74TWiui/ihUsOgqbLeBtvsJUV2+dphDbHMppy4q2fCXn8c3BL7gl9CRhi2950Iv/EF1Q
zsh2eQSbEqYJOKIICVi6aIohkmnNasm+yjIvdBsTqqU0g/5UCKTgfWeMjuu2LjzMyA+mddk/i9zL
AyG2rBJ0giIRQLgZCE5I73tdBmT3ENs+PahMiiWMcHqCIgcUZnTa/mUWNV/jwRS3cZNZqbEtfxld
8dHco6/Qd9/bTc2JpJURnJVhx7yr7r4RfmCcTEy53Klo5AI3pLsj3zGvsjt7TJXQ3siCSyWilxfv
OgFWOsFQ5p5KKoVXFZJdspCFKp3rCkDyMAaHAkG840szIKs9CMtvAEORSNyxUWhINpQ2iftqf33U
2uvIilNjYRIlcmunTepaOiLgz+Z7ildwCMfYlMQw8pone0YXskAgDcwjymBkTPiTeDaQOyJMGTJB
hbm++wSbNA+CbnJD+0V0k45AY5M2I8VxnoLvGpFAnWLt/i2A30mrJDTC6MWYQAjLEWl6adm/c5S/
5WCxfI92O80oIxn6s3RPKRtn3fGfeZuGPltojxN0Ay63aeswyzcm2APGLwpK+uJvEut8yY5Ha8Vi
2ljhQwzQ1+esc04lzlx3AH+h5GWrmvYF0wzeCKvCEqTTpJV0ov/Du6uJvgo31+XAJ6tPzSS2wDp8
DZ4KUczFSIJXRaVuUKRc2mAUNT9aWToCpvvSexhDgBHrRO5g370kXZ+Y1pw+M6snrJFe31cff2FE
VuBlP7II+6H53+Yf0hNB9M/Xg72gGzGI18D1xR5N7EejO/NyzmNenAx6ryEhw8Kf8PtKg9bSzhQm
/spQxxvv5NgLe3ySk28BM91eaak45r5SGwOSadXBbxnKmLx0IV7PEGZ1AwfH2GLouS+ZzGnhEZor
qUQhycMDfralsFNoCatt/56jXZzT5qtF/kf5WcP9zNyts8LckST+PdWx473KWgRfA62XF3btY7LX
Jx2NMbsnhjYVton5JKjSOehecJb68m7Sinx1uXBIbCphLQV51oTMqKXnVBVkMUODT1IqGBA5dt4i
HRrZiJjaOVd0NHcuBQG7sX1l+pg/aSQR31RzHwTJqv/Pb9XuQIvwHp/q80y66eUjlXqt+g7t8eKz
doYqHYO44P21iiowfqiBRtNBw/jERkYwNhibJ0TEJtvBvYVh1qIFMJp6kOv7p7gqfFr3QbFsw5vI
LF0wAWeZde7b1W3mRpp1y6i4MHIZS5sr1tziRgO2T8sfzR2NLcUVEzuctw/2uVsUgzcUra4AdhHz
u0UaNFvM6w+rV3+jUfJRL5z3yrChixeuv+N7uH0ax7YI2nxXiS//CcPLUG0hNtDVRA9jjI2lac21
RXkAOd/Y764x/QuDEOxuYi4Ibw5uZZVbHMVVUq9C1eoXTH0ns4I3TRxoqGtZJrKQc6c5Ni0z2gVs
t2pYAtL3yIEv7cV13xselFsvKnAbE0LuKEHhMn5Bz0amG88G2INOOAR/SQIJgBse/dUqE3IU5BJX
FVYdIcoZtWXBrPIbAW6QOJHMuRy5H4om4z75R301Qgr8kj5/LVmqjMr2tH4uEavuS3F2lWdqsnVj
7OtjKIknqtHoxTDCpn3pasfwnxpXM/gspWr8ljuHO+msf2ydVqn1wlE19/VRZGGRgeg7c9uTB4of
J93fnReMrUqcQQ1dn6tnvlzkYf+hIotBZaJv1fL1aiaF/jWQHweE93L3mE3o/UFUCkhqTPyeKGlM
MDlj/Qspzwa7lyD1naNHMPSWZvE1tbzBuUUbQH+Adx/Kf0CcIXqFqpGWd14XPWluHC0I1d4UZJwe
j4HJFUZllfrJ8UaX47ZKwXfx6z1W1qzk5rK6IKv6NwYKSqGJQHDlPGmpkTqkhYphmpikO3QVHn39
vf9kHavDYhHPzpqhF+vMQb11ZNjLWgIo6/CxdZMV2u2mvNS6PDTP4720rGv0enbeZ70djZfxWZZF
SMW6Pi16F8eTHHeW+uPhMHCgfSzKb6NF/fiT1sMRGGq50F4wtoJMw8idUK9Nojrz96EQ3agtkQ3E
eeh47OksIrJeXwO6mjP1kIE5Kyz48roCfniqW/eZKN94nEiPPMdcewRBzx2FTj+Yr4bk+MeI4U6H
SHEL972OE7lhjUihE2tRJ7vU+37ZZ9rOUEAHIyl22DZt4GajqG5jHkkBlU9NYcdQPB74qRXyTb0W
mqFhI487mDwgrILlJrhVZ87YZ1y06h4EIQsWyDjO2p+VORtNFTHaY4F31tGPNKzApbruR6B0c96M
+THG3Oq/fhhdogTB5Q7dHtZn1wN9x6zcY3NakXBR81bgjXnvUSldlDeeIDZ7PdbyKVrlCLaD703J
15nk8QYfIT9Cm0NDTHEERfvvgQIvU2NQGtD4cL/wmCgr0HSC5wR0D6gDjLk01YS8A5/zeskl414A
jGOQ9cTG5dlmSFDNDCuq69nKnbFtIoscK6hVez2du1domzxlK6zhmoHG1ib+QdpDdFVReOxAg1Wu
1gK2WW/CF0xvCrvNe3MVgHsrGAZBZaQuR+nhWpMlm75T0N0SOUWUHNxoPASewbdIf+Rayh7eOYIz
MKY/ZIGXS0iIF/4XAxR8oECRdiFLUepNkIeyS0xAB3awJXP8vtVcMkg/Tn3HiWFJ3n3hQ36QTknu
UJJUb/19ahnR9p0EmbqBckGty2Cnh6FrQ4rItsMAmn56aBC7n02yEbsGnYtUa6MTI0eXV1u44Rfs
SfLIf7UMBfzz06vVoqj2WKNeXQSEJjPUqSuht6yVgwbFQybhWMy9hC7M2zaf+lMdzvmQ5WMLFtlw
j4J8FMnk74+VATjupCA4TLL+z+ibEdHZhykGdsyCPjH5rMitiAy/ayopnfsP15w50Q8gmRrnxANO
4RKWUFJE+tONnK9iYAReUJn5gP9CXIeStdyTtre7KJp4c81nZYJFh9m0dbeS/y74CKZ3UEBW9/xb
tQ7M52+f+swaEEbOcHtNJTg9HtvIiUU0Dl7l1J5PhHYwFKIbPWF8MiTfu4N9fWCoFw2stdzdukDL
9HKbQhMYPQ0gZcEx/Y+7/IuCgUb8uyJ5EIFr6m/Eb9c5u8KQMhdCiW9ZT2X3tsNTbXeXF7NmjqUl
NTD4IxarclT009kOfEtAn1yu2dgLNix05fyDDNQsPOU2PRgsuZn1LzQSmxkj0vUowmDlvZlzi2Ck
v1wmcIp3kGCvAChHHRHtiwk83j+PK8J16VZUsJwOB9RiIEcQGCcpzXeM8VHgBCtFyxaWaGdwws9X
/TSiTah1oJNx5PbW7d2E/wT52DrBaCce6b0hABXdqgvV64Kr9LIUkVq/IrqzX6x5CDo4R5U/y3J7
dCvZEKBqPToB++Qd2b00jc4ScyqgDu7mm/v0is6spxAg6PaxvsWKsRepSQLyxO5K1eEpxgMmNSIW
5yPpPkSGNF8yfhFURB9IqgAuXmSxBSdAqdccC0pGSFC2D2Urf43AQStLB65ADt3cpG3BVvSPlrZO
ECHQ8mAaYzsvsv414QuVWMym6WbmWUDqD+EIEH/E1V0o6e5gK0hqVGBKk6UonmLHb4aZaZLXS8D8
2/sG9RGdxjSXhKgPNLujGnh/nnbEWq/tEyfB8n1NPtfC93avl1iCeAtaSfSXIbjOLKR9cJ8Quv4b
jb4OR4z0P/7F5kV6TwtwBHKg9aBAMHJTB6cAOa8Ciu5ptHVC4SH86yTvgH1fD4gmUU/pltJVTtj8
64+a5UL9oBGLjV9bgNP9WcFsQ/AWy76tRoc+Z5zzBhbj1Gl7ZljVa9KnwclBDBOQA+rmRsD7ai5b
hXJQ5mZGBM19b9sHnGWDz/Q/qZ1yM7+jKFND9/5kpaXh8WDPKO9Sn5TGa0LylyJlNNS87/FebKi3
jjy4REoZJULmul0hLPERCuQajq1lonWoVdVeBU9ki1/0hA9Q8KrNPKh41lYWK5I+b4fbFPwYDMtn
qtqg9SjbpV00m15GBLcmklK5muR7ScwEtdTL5WHWE0UXSBN3QWqH7E89IqjH2UvsIz0vSd9OJWSR
NoBTOVvWVi5rPcWUNXEa5tqI8D8YEDxkQFUoovNBQjh7uL3v+bA0Knjqnjb8O1lzmOSzOqo/LHtC
6vlfAGeZh+WrPLnAojFYbiOeA1WLurnXcUypjY5es0L9lfGMvAZRMrk4n0JBZcHAt5lJb83dW5L4
cPFNRmSnLIax6Qskq4/6bkt+cCNuSO8q6ZK+WgBk/5LYJ4LYZE9zbJWl6wJFg0XuGAQTDjcxN/mY
uhqhkit71vyNU1A+zrB4k16C+JqW9uE1Ei8k5dQeWhks4ePj/TSiamPSTNG/BUhZEqzulI55j0et
rjbYdfdXhZhXQZsep3KRljaeNlvBmekBGupNh4WtF56Fl0su7VCMb5ZShs2hfESnhw/9j7+b123M
6lqHI0SYKubz5Pz6oVkD7S4dVjR0gw4Ek0kerGcPgueOxhU4zFjAc9Tj1L+FuXoUCDBtnqTRze7y
qpOaakibTHDnO4j4s56LeuOd/h0SRv7g2ooYCPQnRr2iX+YpSqgEJLacjrkWZ+HRowYe66ephtHN
xDIihn/2Tw3aQbuEJkKsuVUMKObEzJe7FCGs8n4QiF3mpIVHAyzVjDDldMtza4ohq48K/V613KNw
qi10wUxNPfAfhUgmL5sTF+033h6oO+Z6EgjFVmrUf0kVk+0qLd1AFDisc9454WHJWm/K1OyXIziF
bNyDKn01z8WBPkUN8IQeHa4AwggbM76V8DaZZhU70cd676C/0aetVo0F6wK8UiSURVW8sSySWPTw
3OOC4scDfhzIdlk7mcL8+pp78jfzS/pDocHoY7WuObbYZmDYawTZAGV2cFnJ9VOCpCCd3k8p/2VF
aVu3xBHHSavSvMlTa3FooWErCGrBwQHWC2a9J8M9qp8QHBAk0dMUPGYwl+qXuwYWwSHQjcDOwMMm
ERCflBJ+3o8rsVtEfmybsznBidRCTQwl1Gy3l9wE8HXO4BZhsSHH7ZOF4kNQwvjWxdEBX0lzecRc
jYq1V7DFraF5VymwgCMydmxwJCTC8wCPAlolXlBzDZ62+rAsN/PB6RZlqMc/cPH1aKOcngzFVKFy
Zf3Uq0fZKOOw5258Jt76L/+tc+VvU8ONeMdhWBRSgb53r+DwKrFThw7rgO57ZpAXpl64s8/hwjum
XSx3YYw/7vbEfUNpUogwmeTEvCgQfbQFDaB8DVSYkoxx0ZE7uWTQtwBD+mQ718TMwS9f6X+JQTyL
4dwYn9f1MQWupey1yLD2PTveMlfFji9kcvCLcxiUa28S95T+y4gVBxvXDcDwAweBHmO0U4NsXHJb
xYADbUskNr8iP1LDS0hweB7ZIz5oGC3On6Iy/Ku31qLswmNAYIo6Q1/sKhDehzlYXeOIb9pJ4UWX
Tg8uXfuM3O7cmzYf08OISGRmIN7CRRYntwRvnJIJ0/elp5tHnuYlBkYw1BZFsjjN9pHsudBQPFfq
EQRRfZHBGr0w0tY6iL4YbpfMG5hb33dQu6rvBQNo8n4PCCsy/jpa7BdGeJlAN4dRLrcjyV1qhGlh
DuCi1YmK5jBDBJK35oQTlZYPmheOTejrIpwyQjRYaCD0muxV9Ftrk3+qjgXwLPf0CfApTEjUW8Bz
FCuFntWfIlu40WGbq+yGMj9YtK33+AsgzDeQF7K6T2M2t1yv1Ar2J6+iot8C7+yPrOiBm2U3xvY0
mqnVO0y7Je4glQKmCggj2go3fN0UzX7natAkWG839/lB9JTd5lKXeaXNv5mQI0jZZjnrTfc3nyVI
2oEN0dm1Dw3Zp7mQy+4noUWu6hCCZ1bQ5dGJYrLDi8/3HUmwnXg2ktuhsXbpVnlGbS6J7QF50JoK
xyLn7hUDpnDBkO2UCWBBrOUG4FjsNIiJblvPkIIomo2JRb9euc+wOyxvTrgJnfFueoae6wH+Mnha
XNP9HQ9vV/JyDlVmRGPTUWKlRhHF0b9Ji5xzczr+MnoALxWt6erluJSMZPNIDjyLSw45XIrBZCuq
zSNcYNp8yaI9ucTtfoJA37LsdPPwWqY0x8OxarzdRtmceW8+ioDCK/uERb4Vw8ypRVlzj1r02Zu5
VQY4CCLn9BKdazvAgSqceAKHbo2yMRuPWD6TITwxGPSGaSB0tG3+onsLKtJuQ2YPi/ApjRPCe3h5
8knX0N1dpdqjOqJF8d3FGoxbQexIDrlDHPq3zYPBAu/aBBK/vYPQSIR+ClVc+4Z2glu7zcVNjrSp
isi4mVZn/0ZMhjyrZIHbwePvgeWTrFo9Ky+aHOD0P5GCP0WO7YVlLjdTfClfaY/lnefA7c4TyfVn
eTAiiIMl6fUcL+L4pQdXqq0oKtV/3W5NV2yLjms2l1GKc7EzRdgRzHKYIVVlFcrdV9NsZKHxEmy0
n1vvubkUoCLFKooraqVW87fIcLZuOefq8AlASil28lJybhzle026xjzADQv+/mQn+D+5s8HbfM7p
h/ujyUrlQcrP6TawyFnPQwd+9SRFl4J0DF0aokYb82yN1GUNhBMci/CDm6m/GSSUyocbH5Ig2jYD
ojyhlLG4lvCD0ZygIX933R252sD+aUvQEhVsDrTi8SQ47s3PrAwTNTIgRRHs/rqWjDz2k6OI8pFw
NlsmHWEAYKrrohHenHX/GIgEuacRazp0uIQNtl7TgoI1UTB1MR2ZfWH8sGgOzdbcHTPjAtX4lImF
LqXsfq9j8UJ9TVO/nPwK0AQDS7ucfoqabGTn534NzYtbzOz513HEwXiqZ9B8maiPWkcS6QjU2fLM
YbEeoGGUXTvp/37rEmct3EOrJk/cEkuRwmTtTk2ZWqUCp/iven9i8GZEVQbHBvL0eVp5Ms0rMkjH
OTio1Ozd6tSGeiVX5hPXDJsp9A19nqCpGFhl4wh37wHMCPIuMU9khk9P7ip14N8zQMSVzOtvQGqM
PnjMXQCX01qDR/DglbJzo2Mir1qIEj2PQPgtANXpzBronSnvKfYHxd/a7te/bhmMzLGxelXElADX
aKsyxoXHoxRBbrFSZ9CZ2qfgojgy/ljH30DK2h6s0rhfKYa31XSfu8JwD25YH8Fs15Go0+TLfKQo
mGJhJTnBe7yCEW0Vt6nmIneD0SUPRXbIJsQFzB7YYChJBWIU5gJ/ZLm2121wPUKu+7cyhkVE08mh
GKaDWnEYcTGzwJ922dqKM8xxWbulS2e6FBls8NUCAqbsVVSH1qihizBIq0Nbz3U2illjJd2uz7AA
NJaIgNhHkDdmTkojJyCxZaJX7vyFmEHKbqILl5JCRNfbHSdNmZKyeNmTYeLtNuXYdAJj6aQhuSEZ
7yPGdvsIngkpZZrOirrCiGkSIVAt0htA49E40qupmrCK4+ShSEhG1IMnWTC6kAiK4CKQHhG0nXm/
5MgrGw4ak4Y4xPR1D2nTcbtDjU1Sk/yF2qbOYfjRHmZjLuvFH/6Q80+9oIEPYuklkaZAhwnFnZ7d
6WUunWms3P281xivlb30QKRbxRwgUmjH7td3uYO3VCiU0MHHYZGw8RAVAR5TPWmo3HaZSwgA8wNB
WkE8IWdRA7nhj9/V931J/RUdrXp4pJmrZFZq9JvFuNTem1d/UvDqOQQZX4JTZub3fTdBWfw5kPUC
DSopRsIxP7YAtVW8yLgZRtSmDkTfuK6LlZ8IpmBr75E9BP8X+y8dAQpxPgI+mAP462Rz/4SpjfEt
6DisKGO67TqZZdJRxLbhfNpVU5CpHDBaGTSzO1m6bHICiipgOmnJjpog58cRf9oaEz/Y6A/Y5lzu
fb//AVVjZAjbYVOoKmA+roZMDn3llRhPFFi+XjsAD8T+pg1OTYY+wLJJ0zo4N8twMUJceQo2RdpW
eeluyZr9BuIxvxr4Xl5XzdEQniK09csvOtPZiEODhi0B+H9DeKc7k5ZiW3/7KDxnB/41O3UD5++t
66y+/IgKjAT0Rj4wmJWRPOsoTG8rGLsuJXW3MFMdHuuBwedSD08qMhLwl6oSPrVtISx6As2gckqk
OYnHnt/5AeV+D+aFQZEStUgxsMQy8g4/zNuFpUuP8xGGj7ZiY07yhbWNSwwPWmCwtUml7bZREOdb
vdSc28198/dFg87pnL11PcYRGUA0bby1z9xIzJXIPOzcGy1hZ6J8A+PYBORrd/fzLT3ItfivF4M5
1FAOI20RKAmk+BUbNtIYNhmd4t83uscW9V+M0sBxA1kS97/D62NAUt3kgAPRD8LkS3Hs3j+xq9W0
pF6xSU/e19JwXs+X1UeXtTb3zZ63IWf1akXkU2z80jfo3Nk+OTkSkV7LmCchvpTovC+lvPuP5Vui
yWh6nB/hq/0U9F0lBkUCRTlWC/YtDN2eiMWHxLtxRaCVsaVvMwk8Iy2S5eJ+kEbFj99rJsxDudAB
9r1+zqVUYaewZ0otwzH0426KP9ZTN/dfBSPz79ysILUIpgRCry8ZehXpAXOgmyCE25ArQ4ZgjHFK
Q+s3bH2du6WAoAIj6AoV4jALoKbK3EeB+DSDrvvxq7Vkf1JouNxFAhVSknkjjwNRGco1bMN01hBT
B0n5Y71NHB5mGQ37YLQeWNTyfRWz65PDZn8gOFkkXJWoedCJtZ1asyvSqYwcAVPUSvqxI89FOh3Q
TAEr1d5sFlmr8dh5L5F7SoDVYbbAu3BQhftmbLBDhbz4bmTbKV5e4C6hqk/SEUDK867X3asbSKN/
o9CRaPMw4eB1gsHCOAir99akfSAgPsY2UAkPuDehkH9wslDggbGPl3HUIhQCZDDkzS+LQ6dyWbzQ
t8TQDBG0W5Ee/EhsVcpatlbezLtTPLyFdemrgfG2On7o83ZhYOuyW6ijtA17ORnmQhg3xns1yR2Z
M3uu5mdnEJU1P4avmjpOXraGomiQvzBlgZOSijuPFNXwF7laMW/iHNYV9ZuQuIuReKx78bpcFigO
CmZzCPDpkLEQe3cFFfQ33X0AlWgOutPU8EBx1PG4PNb3rSn8ucfhOTvZl1iIvmbZUQCRneoysM0t
2H+umDizdHBMCu8vmCgghCy0XyyNi0lyUo3k7reFDwbW9V6VIU2JQfaHA/j0mE69jtm4MDdYDLtj
V+nBbeHFTueci7tl4Lt7+vsqK9Uq2zVwtgTm7OIWSjIh3awXue/BD00+2JdrNifct8MZptVjmsmC
zTZytpwcIajMwtoKp0OR9WsVVr7xvCSsn4Jl1HWd4+NzyJlHYWYE+d8kQ9KMemqlp5YtMvpKpu9J
aPZox1ZfBSv5STMIA3JGuBgEUiTDcWzljGGPQp0CIiqgfd2uxqQLA/ES9fcAutUTL2SNRsan5miS
Aa3UoWTURvvlFGxcgF9cbtNGCdKQjkmGthKWAjVBh6jxQ7N02LADBiT1w8DkEtD4up7xlaSlKa6X
5shcwOtlAYj1J/dcPCbadtFTWgIaULeFQegy6aoM7Dxz0qZW/ulK4MOuEClxX+w9ZO9Oze+ziX/N
Mln+cUCR3d1IL1ioO+AOhBhbnhczqrrfn6hdUpedSLPETrneJYaKQlFOnVy8E4Wry4pdv2PeRU9f
qexawPbKCyH3gd41fIGP7HfohT8LCM6wICH9vbeZzJgp1sGSYEa6/QWUFlKnvLOt4jSBmlR84lqy
Rh4UW5MAWte6zWS+bPRLe4kjTicadOo0OfsXBnJ6Mf66dL9xaQ64UJCb+rewNPhhb18Cc+G43fJo
hS1yZrlyu3j66yF3POVePe3w0aLHxV5nA6RoxsbYNG0HpdwDTQ0vEIz0iBDDxqa8TPTkkeEvWKqk
6JfF8dNToEsKyY7EBIApP4Rp7e8joW+CZ+MdqpLdI0LAEQBMsVeXLeBcYhygdPQZxHFEBOY4e3yR
KCKXcOCjxdd0I3FSBRo9h2dl52DOUebGYdnTVeOxlvWo8bRd0FxIjCj4K8XukTQ66vSNcq2slKJe
0Vr1qvqLpw7PV6Kpj8YQjkAvwSC/qwjGonyO90irvclcrvoPbMcpV2BfB18btTUB8rmIiv0UWrFl
b/QxRCNdkPlwsBdU4wwb0WWbzTQIveOtOrosj5iuMLmpA5gq2w/7b583VAmUAbR3IvWB1H7nf1XZ
AdQdF+UBub1ucr/6wLfD8jl6GcfYmc7O1uaF8NZ/OJKZDU0fIdyNBVZhGP+yXx8kVzUFt7BCm1A2
PcHDOgfO2Qd8NTp6D69k3Lr1EvVgC6XRkyiL9+bmB2jdyqZf6MejAcv7HvYwdjtsLg8sXYdd6md5
uoowKoxnNo3nx5aOg0j3At+c8mnXDV3x6wyyTUK/+HmcDxdAaQpqcnAgC+iVVS/Sgc6F7xZ/z1gG
m579ubIDSoimNMB9UZ4HnWQGL4xsAc3RFzsFVZVa82T13SdGPEkGTZn65G/+QQPClDojUJxGLlYV
TpeTodebQ4VvzmAzp/JVdPnAIz76pOoMrThXD/EJCTMTj+Clk+FV8ySW1mVbM1XGVm5s2E4VHI43
EDUoui5622xqPi7qH44hCMML1IfJrYwiwAL/8Y/EpBkE+2hdFwktNcu1SRZPhp8Pb6iWrlOrBINP
dLguZ7ocNGmErSuLtxx77MEI6hHQZ5oT19hE22gY2d85ILroX/RK50p3pmNBXtyqF5Z1bra5YozX
yo9sb/bRRNf3NxVHUlFV7tyD21N2BGFAALEKKHjsdM/i+AO5/xJN0mKGzM4E7iBvVddIqgcWoAf7
mQGhH/l+56zQOlPyBZArtGNVjlO/XNu648+HUdtJsNOZioD9wpo4iu750ZQJ/H10xmla/rwqp0Q2
8GFSRqHJwpE+Ptn+cBTRi5Au/mVsw5ivlcDPJ7js44J9rVDrlIk/h+8Vh6U+4Av2G3un8tgNBdLy
qkpYCjFXlp7j5brwO4S3R4l7J26mFMyWnGoqBcQBSZKrouy8I1eeTytktD2FO/7tKzj5Wl3k9hdO
YEBv5aA21m6Vhlp6Y1FGbXs6smWhvIMqRPjKO5lS81B1bMBB3450dPVd0RogsMmrJ1J6BMQTvXIK
yDhZglOYPzSpNriQzS7/8xbP9EhsEItrjqpdnLeBdiEuVpkxlNibE1XIhEeTVNw40J+gwux6tUvL
0ZIXhdfHBAh6fct6dIIVInz66KaD9cx9+5TUzd7kLLKVpZMsrUOkUQH+2R9+1r6XEZR/AHa5eLvS
fpDYbkOWCJh5DNvCaw+qki1D7nGU0CgJN9jL1bLp3dFiz77GJaNQY1CRPsshVLtwB4mvz0XJh010
KRCYDKzsLcA3vNHEiaxTh6KQHjqSY9lZS/B6KlZ3xGBVAVm0LYd07WTcD0fsnaQ7S/TrEoc0gOfx
l0CyaVqJI6oLh6OhFzzpYGeFOoiuXlLuqKrM9OC0I0O60+IE7173YrUT//2PecX1TNVQCkvCsh2O
Ixr8Jky/9go75MkGjGHshD84lngGV728K/etLT/UQp6iiGp8Y+8N/MSDhS2rdMlB8B7XTlulo+US
BYHgjLcGIxxw+BB1BCCyzj3V6DHaL8QYzzJJaHdLDEmeYtUHdqcF0uK0RqTGKb/zEZB7Z9MYr8Pw
vDo+EY1r0nBuac41G3/BnVpkTK5JjxeC1dG/Y4SWgZUifgnMPGmrGlMEvUxhDG8gIGPwOv5ycNjt
yjKpbexUxvMCFAaG4RvZzHDEGHljYwYO/kmSZ2hUQu48yQTdcMAVUvD463sjizdCCCtXr9Q49OBC
/HgGmg70lIXk1iqQFtFSDCoxjS5pss7ajFjvBy7kkzNTX3w52BfUIWg2+w/5SL5DISTN1hy38DBl
HUrCRvwtFAzdez1/2am07NozDfU+VZdPaZZu3YiWP1N8GulP9SMSfek1fSZm0u61vBq81UCryy4J
w8YYfC/EqxdY067MlqlrKHPh0urku8MqugKu5cBOiDODg8jv5hlK0tHeI51LlL76uJkG2y9xzf8L
2rqzdyGjzeXA8sneSxhxeDhBCrlrjNzjhnVOOykQNnscXLkt9nSE90ZqW508z5KZXViBkTY/t34F
+CJ8VZKWLTsiefnmTy16YtAT6JaxnAeK3JMLYq8kU8I9dlAlxE2ptqTH+fIX3f4apgd6LD5ajUzN
ZrbT1L5X/lmropTgGXksXObwxTrfz67hNR8gb0vVsO8olZYqm2XMetpqqzSr1xK9O//yxNN8Kgnp
i9CTYVdDhfZOXClO4ynReqrEBdxa+XvIW/J7GAdJfAIeAL+ywVl8Dj2GQnx8enO+bFEh5/nICoj/
cOgVPcpwrm2TZ70cYW+q57XUuXOZ87pSYgGQ5cc373Fi6dLuBeXXq/RmTucU/pwFj2n7NtmTfXZa
EDNqT+JtdfbuRy7wSEjXoaySZNQMC5y55wWtK3ic6UMp4DTCtMrgV7u4slMP2/zDXRTNaQ2w2goq
YrJaU1mxst/fH+jib+juB1D0e6GgIsn1EVPfiR3Yu3O48vmKAwxkv1CGsrTJpT2vBOMz4iEF14uX
5gLs0IuE2sHK1Wn5b5TqIPnKrKkKCIhs+5dU/kb25FRx85TUXp9/lQAg/t/divGoFNMzZvkO/w6Z
PjuLF+hCitN38xD4PFA+uLOlptZdq6MX4vl7/IqTAm3jq3W56Q+WDtPqQHziHiUJzUHTkftiycsi
NQ4rndzDSwbu+xWAXXgNFWjxU1NpxnSUJ+wiO73D27sAvHroazk81NFauubtvvWHUF1NQlzTy969
C8tlJpDSRl6DjoYjH4WDbxQyoAEK1uygUnG0WSaW//6O+hcRNVVWKaNZ2dcMSu3vNYdlnxLfGVnX
TOcOUvtcDivvb5pinPu7BzmBnI92w83rBnp+rX0evDIjjK/npp8X41+ZgEq0GuINREDfgDwVJJ7F
Bitdj7q6B69GokRuhgDnKHrlWiFjfSHO72NhYQxnT6PpCCqZjuYpMFY7/c8gh0hQdDKXeNTp7o25
fR396pNlCT9EdED257Z4vAsSfErNTxUMyBkvGLRpA8jrIWhxpXur8U5HNDUdpCS3NotzgsZMNqeD
Xd305I17vn9AZsbudhMG5nkvadHLKrSJBOhFKcMZp7XnJ0xoluc+2wqd8fXbF2x8jV1F4SN25FQd
ISeArN2ibf1evvt/h3dlnIMJK42UAVcENVVpEiF0zUwz8TU9pOrrzwG7KNKFFsz9xz3bRMwvJdZx
wnJx/3fdoHlv/BYh/DleLQxVl3iPnTUT4W38nykf0FUl9Sq7RCVszBn18ThJ6pLuUFXfxSpx7kRf
txx+ZR5K12L9wgbBO37xI8pv56zIMu4IipVgOI5NvSCS3jfDae+GOtOOi36GLbb4Szq/7sE6eVxL
XaOdraq1AdsXt6dKNUmkIx/Ehdlv/z6Mw98dz133JQ/9Am+Xko4YiPXtBdQj/kVrbcCSEe+Le/wV
ykZD+r61hFH6ok5pZTVRUgq7oCDItnJPiI5Den/LKDb48iRfzwbCCX0asVxvrFKbOBmL1LPmZJAZ
L7fIXtmKL6JXyX1KMU3t7CjGos/JHzVD98gkXHEQ02cVsOl5fqZTWPztNXVJU4CpiwqwDEglSUPe
t8K+6z62Zd5rv2LP1ng+cljP8FPuHYazkXlOPl+YiB6KLvTmwzv40CTSLpqQSZZaZgDoXmuEU7wQ
GEbJo+phUTII2YlavcD9+cywUChfPANHkpO71jYnoFHw0xbMJuARm8GoqYFlBvo5ec229dhaHenc
dQcdgJq0laQr2JucwnnBmmUAS4m/6oLMPng+rweLiREaElSiYlBOuTKIL8KDF+QsP2XE8v3BdJeb
X7P3uArhwvsKuVrcRzXiYyBUe4l5MbE9DfdQG4q77+EY4YIfYAb0Aw0B5FonZQXCbELHIpZP8Yen
WSDfAJFfn9N+O2OS52y/zY21f0hX00sleVlDlL/vo0TCXwkq9NQJQOqo8tr2Zg1X/k6iA+eh9IyM
PMVwj7ogOBrL5nuZA06fTN/ENkilNVVo09PytuH74MjJpY3ywbG0b+f0h2jNqI/2QnJRU2xXxwm4
5Hjh2J7dxK6FG0Ug0EbwStR6C4aHG6hgWLgEczhLRvY4nF5ClWtJhxJB3ijJ5ya1/c4mBVu3UyFF
phYvjFY5pR1dpavuui5XtGy6F3ZSfOC214WeNa2nWFaQV6SB2bRiVG4VCQHOmDwNOZX+4zqdEXC/
ZUwDy4Nk3Rz+kRmup3oLk6d4m1B4Omlmr+WQsSMmhAE1pzX4zyUFCW2evcdBANgFxBnUp7JVKT2y
S2vy+t/SMx8IlxjV9/ov1oWGbbnPUs87lLUYjViunK6xjOsj4KYbGb2ft+dR8LoS7pcOyEeNA98l
WGXcQdp1KI+fhChTm1dkHX1OaiW245OH3Nf3wV/NUObWZbAp1tUCVVEPa6BA4Fmw7y4eoLX1JxaA
xVDwRYKeVY475HSTBNEpPGhLst7Ea4E+OXMbx++PSZdXRrNfFUBFSvJpu0nofJK1XrcK77caR4/A
V38iUp0OzMRvWZhI0/HF081S2IBHyXZincFI26SlPt7ru7LteFqkDe/Af4zO6dyBOf0Ozpuy/Ko4
c8PUQu5NBRkNO8fJsxSJBX8gqRHbsGAyuaKiiruYKWw76J/al8FEYgylghOouQ7NUHClPjPprvSw
t2bWT00R1Rh4WjVbCWp6gKXyJwdjqjaiw1+5kXPSHTM//ylFsrTB3/mkgdUDBRo7kbamGmeUUg3n
6fYfnr3mwnFq8ZN79J6yKQoz3+9RSz+xmIStdh4CZwe+XObCx0C2BflqWORpLI/INfbNa2DGiT5m
LalE2TiuKCt4jzAVz4gQw1o26panXua48hNpsMfWxt1IxZnrhH8O++7MTLFl9gLvPeo06j1UIKzE
kb3wo97aU6iNdpdefTpqmXjYXHreaAIw8c9XvkuptYN2KXYyG+whLDY9SZe4cfr3LBl6TnlXJWTY
e5nTAGQ0Mj8DilBSM7wJQs8isNGY3i+SLthy6sc49P1she52uzzP/ZhPBGZXT86G/JY8oDEUsreR
hJ8AgunBa9X74F+pxafmBPj3WXX0KBVPxoqDGrPTDR+fEY9dp4QCQFYXJRwvBaERxBaU7ARpJnaH
lYv0T9Gi+hxdXKVwcWcqVNbw04BAr1KWFf7aSPQODz2UXvZzL51oHkomgGhRKXc1TsRrWbkSLA1j
C8dN3XgZyo9NSpwE8lO3gsSNmA3i2zw0W3TGE1PVgEzexpm+mMUOIhqTEgNFlrcD+iKvnYDYWLrm
AcK1bcA1f//mrwqPKa1RiDO1P/KhdD9G7PYxMS32UtxNTRnSIVP0v/qvrb1G/+LYh9R9AtawHZdj
/iIovleWrzUji2j5lM615KyELa6tFMlCfHI9icEyvI2mAb1TtlonNNd1fRPgxS1+Xad9QLfPZhmq
pLIgu+6+I5Q4HYX9eYjVcVfNAflHN4ZtnXHFxdmfbrs+Ds5gQhkeqQsoD9VhQJwerCpZFdjblIid
3AYmKxlaw3DgrYDxLsmuSgz+OIFri5LNVZat9n4b6I3KaufEW8ID3ws2mvAdEXXN5XJu5SzAhc1f
N3eXuDbQpKbso6mIu4oliHToKC+Vi9bPLzwyKDc0+cEDMpCWnlZnPtO1qJYbqBFiajbOxoDXSRPa
1olasq7y6vlQJPI20xcaDRHBOSC1EZaqtMngmPFUy6dbESD3bocLuIGJ7McIzvzwitwFJdJzqNFN
Y1xUjf6ZoAfmzmUru7s9TuUJ4zi31oSkKWMr+jDrOf9UpXxdRozl/uQg9pdWgy0Su/d8nVh4Q7PF
L+ddmQkLRqYCgTvHUexv/b/OkJFUUove7d41jjEyS04aeJy5qhwk7/phI6eoG3naE5iyeLLVRiv5
jUoTiHrmG/PM33+F2X3WQ9C9Luyu5gIlSbegOW4xz7NWt0eE/94N53tqAkrkoXFtEwWdXpI4tXYj
oQiOXSGt7XxtZqMlR8I90LlCc+jxiFjcJvODnntRGF5QcDAvJz/b7Z5pwBB/gak2St+0StY96hgE
Mz8nb/SmgxCeA5ChfkRfEWx9xF53ikjijsgHjQqf+Lhkwnixs4K1un74Tq53Mw3DdbTwGL703Gqm
RecnfRkdG05in01KBF5sUHhNpUCda+bGCgCbsXi6qWTkryhkAHEdmUJjcSKaRbsAHa0nnOKpUpYX
eCVe/wQUh6GqtF91Dzp3cP1qksFZ0d5dVK9vgJY2QHBNVaMj13hjyZfnzfabCcjw9CQNKgW+SGQT
5A5NwGS9Mjxu71dCNIKyDOK1L2qOLEt+6IHje9JYZOrnmouRc2p+PYyE05HIL85Z5dB6iZ4g9W2O
Ig1k2l9MIfNv0xn2x5eaw0us4lzJ7MqfURL+qhDCe4bfCxzvCxN9hOyc8BbZgrFdu1fW2SodBLcO
bFFPcbAYacTAEfEfGBb/cvHzN8F4cs6tiHZ0hf9wx/aWSnZNG+PB60JxwZRNTayqKlU1HYyQiLah
teHJ7jviVT3XDxUKasa49J3cRipfpftHttyBSEVGRopvu+YZ31bm4KYKW+1NLt9R/mshagz3vDeq
aVN3KdGEmIPqKhQ/ZA8D0fdRsMDDMZiD7DLP50j1kwoBFZbhNDiCswuLfGBWorMKJJaS/p6eED+w
DjbftsVSvG8fIUX2vFUY937vgCNDjMBZoUry5L1bTmlFyx7Wysxj929LI3enGa/YxnDAsqdYwHsE
RkUAZiIcxjzWb+L1zj+ZOPdzbVHhH1kGyPvl99lnvbp5K6MkQm6Lru785Q7pHwWbBm3sMjrVBxdW
wlftlorpcvj2D/BAJsf8qo9nl/nER99794nFOGROIGeL/TxsGhu0ilWUgfY+UukZhbx7OwVz9bgH
TEgFmRfrf5HlCLSnnbJMQGa7FDa43zjunaTWynoflng3u9gclLpZD2PMXuKOptACqYIZW/XMhYQ0
vnGdTpp1Rl7m//BLRLcMKqkgL/thFasGgiKDV7zmyEXn47uStrWKgacir3m+1gkeBpf54EYLuOrG
foALyOLODAXMfqMfGwHCWmD6dx1LhKad6KXLPen9nZC+d1aXU5nbBX0R4JxBr45AwXdha0siBR2k
U542MGxk3cUIXHB7dnpU+QrEKY8tKLRJCqfMK//GHy6weHIGERuOAeHDxyOWGTN1el2xvMB3sANG
/1A20tfm6N3omhXYE7f/0AgxBoxqrgMzo+wGWbmOJXX7N08eVIm06UAoxwoCVlUgCnR4hoGYLvjE
TKIkQ5gSQtZGnkhPjxEmtaZKIdZ2DXWRIk/TNXE7XwJu+qd4bQtlh2lLGmWluzl4pTiALB2bMHo5
zaWpED43kFIDP5iZAGyD8+L+slg96H/M4YfxUZ3ueKI8hxeYw9PTIt5uCDeJMn2sMedZr4NFo9Uw
6nIZPgQGHVRaxwtw86iFwTOVUcIOMDPYl4eNrBFLCtwmGaCLW6y6C+d05COp27reGEkU34gfNl+4
0v9nz3CRIrPjVgXJqIC6xzYqRe/wOSB9dLuK1+Naaaq4nYYKmt7VjRU64VJFLda68f3lO9zVu+yC
gGIqjqWFkpuxzIOx4qOzwg7ktaIBn5tdomfpdiUa+qHgeKOrzuXNrNtfjDhHoiawzvmnHYm1aYGm
G/d+zuUbWCZ/bgwjwGxpa3ge2sMX8khGU7yP2HJmjuia36JzCR0MmniiHZ9MbLE9SBnfM/b67ooQ
1m4ohBwlaONqJtVG+YbJvza4RXfES+Hpa5fkY90SHAaqse3kxZl8UJdB6/gJWtEioMzbimmCdqD0
F+AGplPlRnkEeutRpxTTAS9vZ/BQUr55HYXY68NVypeumYPm50YbRw34VYa2lCvZXL2QtEFIo0Rf
Xbut4wAy5l3kNjeG3IP4cl/p7wKep9Xoq/p61NmLEIIltRS0Edrn7skri713ecXlsXeGQgzeLych
T09eofpfFsXh/oMUn8KIUT4iZKnfP7ECqZat62xk3edsZ3LAX3/p7xJRIc9U2CC4ULs9lZpCETby
BcNPbkazZbB5bHoIolw/jtIjxP3Knj6xXnK0RBSfGm8LUGfEkfHi/16fmOw+dGJ1eddIT7TOYNgA
XxoIH9Sv0c4TabeYgdJ4ur3AY++TcXp5KcOo9dTkqtuyuyp4zRkaObiIJ0yzxg8VKUGXmYEWGWlC
X3lzzY8fegTAEica6e4LWBjnPsrMvnpzpUV4Wl/1HVy4PpPRuwyGbtwzkFHYJbwh6nyWyYMNDegf
t5AVWyiiiD5fR2PuBvhVH/BRpqM/J7r5B/YFbqmajLuG9VzYmp9ldQOTDjM5AEC++oZ98tUpgAh2
zbiSuRgqjoJN93d1lmE0628S1KX012853r2+62Yg1bda3mWBArlhCMRIURp0oVq76972SYYdNa+g
f550yNPf5ZYWaQ/mW75kQ++Yjt1zy//tgite4s8Zxdx9YjSNKTOjKi5rkUFsOJlCyZf9eEeKGQls
wmI52Q+cISgnd/+0Xa5jy8lqtvJJbl7tkZ0aPb9ERcFa0zZPW0Qb2SIABByleSULyxefHpZWYud5
q+VRUdUKuFpUYLmYLnzIsCpQwXplWhRCK4UeIADiW0PUB/T1DYmiTht5r7sFfpyaJb4JcfuypyYC
OUlyanNZPMBk+jkJuau9aX6E8x+LXHXfKetjUARoG9i2PloA4qlzIb7OA0Wvf2otiP+iYpMzwE2Y
kRnfTXyVX3P4M1VVS+7jfEypB3K8Dhdd9k4XBTUx2Nw/2yxRqnRRaEmsxuNwYFmGhPabvwchCs1a
Ndc59fwWldOU4O9mmJcYMhSSAQ+iKurHqRZLZAFHXDcB4WFf8Bk5guIWy9rouw9XdZkOwwv2snHS
+urp/BYq9aCxcu53D0QegN4qFmautm+FC9UaM71YGUyZO2qtgA+mzeSV7unIncZhnYU8FDVu5q04
yhngu4lApZ7cpXvR1qpYbU0THOh1XEoZKT2TD27VKwcaoGmxHlo8SbTT6VpMQesKvVizHzJqFjsT
4VcPXLXn/gkhVy4b5H5UqbyVHUfDrnWxQyZk2kbE1qS3AJt+4uHi+Lb4kxo66JyQF/gkY0Hxq40Y
AJxDfbluPZNphdcHRkjapbr5UHdUR0bs/Azw7MeSWBfeIM/Vd3p1boQUcXcPGsh7V8pP7ASlIHna
Re64wN/7y0txWZ/8p0/uINKIggAJlGwPP4bgSuKgUyndJ76oP6FZlD9Pk+l0jm0PitBnMAOKuQJq
ka8zdBbN0Jn+tvMXMFNDVcn8j9atsmliAP0ygjB1gHE+JryVUgNmY4as3Rl1m2uyyFUsEiw1qxDs
dhAOP7cSF7K3nB1DrW1jV14+tcoRcfbvn0t3SFZrvIP33eIL4W/wzSvZb+0vzoKsCPS/zA30nlL5
ko60XyYKxpyVTbH4PRB1MOQk4bWefV5Svt/0ud3Mf+kezt7fyRLLNvnA8OrOahOBvkRUpwU/TWlj
8pLsgFtxquBUoWZJgh+KLg3sDFJSqX53TMD9X7E4fJeNCMohg+ObfUd7Fjtta1XaolR7ooYmvPmI
norVglfbPzqaPlJO1Q3NiWUxvgRgpOkT213D3GaopxLoZUikdIMMQ6Fb9l2kyHYEBBLZcbySN8up
RJYQtWk/zpS5kVCfCBUxCawDN0XLWWdZcEuUtqtBMKjf5eEPOX/aPA2wW5bdcukOnsdJYrWQxeh7
P2hBS8WAIz+KEtMPDOS+Sg47fCdjZjthwhoDnMoA2ZVS/QQDmtH2NHcEceChHttbeaF1wIAhIjga
oCuXdBRM3ggz72WX69vEAPVXhac5v9UwTEOXejR0Mi6ziiXWWDd1pMeTexYlaVoQ4tymH+f36QR0
LuY2S1JLu95WiTMQ3835Mi39n+/QIcPPmXflkaQFHGHEzw+r9a09x9AQpQzWtBNZPDLGGhsOiQRW
h5xXJln6yr56Q8LVYo6XyEwa3okvxU76dgZ5xLK1AAJiaz6n0MmT1DmpA9ZJkEpGf8ixkk/tzhl+
+4PWa0TBrS4HJ4/9LaW8DJ33PCQp9F7P9cWGNT9BVpJnEWJPa6faQejTB6f1Qnr2MKBRevjLnO/+
WtY6eeNX4upGi8Ahk5cljVksiL9k4ozDo/yvBfqBoPcnfsyCG5iQ1xQdCqEOZBwOoc8Q3epL4113
mRwXf7DBp5gJ+WLF0CNCNf1M1+4QRgrSrmfROBHptyHQmS8MtIwnVZ8sNUlx1Nu0EwqUPCu2acKs
H97frJP2qe9+A3mwsz5QmMGe6BzlZDWgUNvBs1jbbtg/4Mjb1Jin5fZU8bAPI2LftD42LkHJhTXh
tH9ZfICAfadQubgULmuzV2BQE504FKOYJ2lCbl2vyIK3CcxBoD8+hoRRiPY1DRZFF9i4o+1Bp9+F
DEQ3LLCs4yFN2tRCtyovO5jxcxN1rPrxoXXcXeGqF4H9Ya3s0zHVc68cKZ2CRZ1t6HFeJE4Emtcv
y5WvVxR+qp85odVLpeX2n5Bbym8Gw4xeofxReFvC/ByMH6L9q/JMoA7yx4nLaKTF9gTUIxKO+LCB
m1YxESKyvupblfjE/Es4tEhhpXO6HJAENbRGdprqNwweH8ujfgLoHD2qhqoVJ1HhFlCutUCnOZPO
7k3gXmcOHE9qog7RUhVx8RBDbmgbL8KEfRDOHmtjcOkfoeG7LylrPNzf0xRK+sIZNSu8fTADin6/
YU8bUrcXq5IM3AIRWCsaeOYICQruPqOhZWRB4FW196x4498NklFVw8AWr2TPLaxyTVm+r9t0rTn/
33GqiG7MfkTtIsp8zTBrcQk1CHHhe1hBj/wZj5C7X3HvlV8XaHvvXfbkHqvl/Gq9rGYAqeDFTZM7
wCBsQ5Hry/W4aw7N5J8xh3I4ZrFI2UGnboOxN7HlfD48a7B5Z5UUlBKNlvvfif9+NPeKVn1sC572
cyaDUKtJPZISJIr6yI3XVcNYlC0u8O7T581xOHPyw/UGGRAE2n9QZKHB1MBOEcICsxTzE6vOrCiz
hh2XTj/rWHeRhIUtxcFUDWjBCA9+0ZDjrerxZxx1eIZd001fVuQO7YcbsnTbnznAQdwseUqYbNEl
JAMSiJ031p5Oz8FaMrl6V9pyQ0pJLlJwbaULoAgouBo4NsX7w/pPSKwVQTSAzkykHqzjoPlhhV5X
Ee7xn6RepLfAiEwunh861s3AdmWrB+f5MvSmEzYuayjFEKrTlpk+1vvQILTEKII/QCFoA5+82Anx
H1pKNw4wD6cu3yTBCjWHVcpzdNaLMNVDqjkdKQoToS8mxjhebQFn6F6vkSq0ZH0Ip9qSWV/SBtXZ
33A0kdgT9rscoV4USQYG10Q26xUXxHK05cPmdXuWfKsmykGLxUy1jD6Bor3cE5MWoTuupGW+2iyp
GC2d2i+STRxhjH5p/xcHXJ4aMIsOskwIqpLxSuRodmISCrm/UFY7QC8VFcl4gKzRHmxNdjbZv6Wl
6Feh8rpa/Bzl8rAKt/sND4mna4kwWEmEVQJ7KPFg6u4j4FFFwyXg9VcIhevnTto3CamjrUG5o7Qs
2bo2W2XtWFd00YxjOgei7RCvFIloWwnTNOcoCyAAGL/aQjJz4DuFuGxP9a3FVOl9Vlt6EztX+gZf
9J5V869ea27rCPEAyKoNg9VDb+RYJEvU9aHVyuTjNgqptbDhILYLato0LxRCtLjPP1dNWcD5uyQE
vzAGgdP7zRXX9oPeBKxOguqIjDuvuOVcPH7evFiPz6RWE32j92eavrxQilVn1IkMLTim5H/w7bWe
fBAtk3CdllOP6II+OJ5neW4emLp6hOMl8gc22u6fvy6p28TAcAtMY0KXDz3htkmB2ybNwaAFUslu
tVSzCAKbkY57r4ZRChoNlZ9JTNYxE6gZAjfZSw2/cK/60SLIj6Y8PLbgeCIbhrITrVs6xT7pO7M0
1k8Hk4knvb64NJ+uoHr6Knypoe0TxOOspTfXW5bD3HEsbmYjLmvJgEk2kK2e+/4V/4w9Mk+FePhw
ecznHeiI2dE8J8+HqqC5O+b9zelH0Dj6CzUo9fPTa3FzdeLCajAC7PjiN+F8X3NvXEZZIr5ceTqM
2E+ZkJHveqwe/C+bZPLatCgAMsCuCLR+FGjyCVgktc8TBcTy5VNt7n6s3eQwtNJi3JIViotIvqXj
tkJCzHXWdoueYA45/naxRO8lj53dQyoqA9cHz26g6mamONtpwv5yy60n+hIStvWZkX4shV6bIc+V
LDCBWj6dpJ0Bq78VXEKLNMTJ5Ak4l9t+4O2o8+n2O7XasyPksPjhom1YsHC7CYVRVtR0DJ9+nzJE
eUl5JtF6vC+Xsy7c0ohsF1cLQpVFNVkMrgqERI/y44nIBCBWN3SYCKDhQI/aSf/lz9V0X1Hsy8j0
wYf1dqM5dnnxNJckjq5LX5SzfoYyH4TrN2B74TksELucXFqDDHdovbs7MKpf4xm8h0Kbqo2d2bk0
pP5Vu6JxRIvPvg6FQzgs7/Db2rhfoG68Rai2wqe21lts0tI8Z6VNChT6ST26Cusj/h8pDJjCjTyR
tL0nJ00QNmRUyrlXfHocDP5O577zdvSB4JnfcSexlz99Bn3/pEw6xAT7ktvir9AJ3HaW4KQYEYfm
J5byBLjGCWLnURUE//5T9BgttN2urG8sIu7XcywuzG2yZy0F2Yx4eR41keheQYE3Qwx0JJ05IQBS
YZ4X8a1wpRDpqf3fVCxOOLQJl27WcqJlvjNxvP1RL6T7qprE4N2/mlUA3FK4289TJSbkQLynR6rv
gz9462+PPUBhqUC34XzSnjqs2AFP6j2rVhBwQliqT2GSQsL9XQja595BEd85w/LH16e0dYH2ybuu
CEEcqb9QNAc++XIvXXrMh9BNeQZj3pLQ5j5FYi8j/Fzz+OaxP3d1+mMS9Ps49Wvv4om4VONXC+X0
MJL4xNUaeHhhUjKNt7yhdAsT3wVoCDOG7xWDVllSd/j+OZ2XxKgokQg68AYAa/w4Nj+wlR6ehbdH
R/5TvEoUoy3YXL09SYFRdr5CRS7cXg0Jv+OmOkMe9I8oqHuy4SR2lsxXxqz5IDYETaXuGdDHP44U
0oZboo4PVa45SozbLAoyo0tnkXpzmt3nme1qfZgrextlZQcaI5UnF48f5d1TbOXHtepHZ5n4FnHY
Rlxk1ilrbBAaXmNwDXJ2NYys8w7zX3nrujlxwWStFtQbi68l2E5DEUtaTTcD7Bo40toH/CFVlbnR
K90b8vMTkICXFau2Cg8vRr1jP8XMqoswO3ijxeA74n7D+8700NKZ1YH59tLkGRCG/TGNsDCOBO1Q
kJl9OhfRJs7a9kUvxllNx6DNzZurxb6t4dXdPlg02sFGoxk2w8ZupjaJjR3y4Cwo1WxcrAnOKA2Z
yMnlwO3opne2zlbdlbX5iQKhAS39XmBDPFie66j3qYXpYdztBLu7i+r6h/oerFuZGyhnxF784fI/
zB0GYEupis+LnmHQ6DDV0gkWx4KhoaGIOqCGYedd87hwfyJ326oObDhpmAOdj6c5/jL/NWwbRxIk
ppKGKxQgNWiSVu9FPZYWoDe+q4jXv5bAkGwZ+PTawGEFbZg6dzH5V/jGxoXzWjs5ctXz8GVxMjdS
OzVSTtPZIULHxZ3nuCXdI6DrtQap6mXXK2PYsXfa+aTTPUT1eM2TYb3EzIqdGzD47OF5hHuWFr8B
ALU7L4NWf/zjztCZJKy4/WLOtAiBTXe+RYf1f61pIPRIFc5HBJoPjU0EbeW1YaKjvZXES5460ZlJ
QymX/htMAFfk+26bNJdlKSZqRRvWehABtC2C4nKsC0y/k1RbyZG4iBHgR4BsO65MnERv09DFwjQK
dftlhoP+OvufZ9TQwE/5ZH1FJySg0f2jjocjwyimbYT8xt2UIISyJ5FXJdbotIsl7xH/lPF89d6K
fUkcbhUYmRX8zvOGXxJ5CW/cwFbIdIHacVIz3qpDoE4TFCVHiH3F56lKAc/HsOsdFnfbUeUE5+pK
8+6QnFqQiLmFKv+3GyW4YLtYG8ljasQE0is+8QqA57mAMm9TRfi3T6+H1dDWg/FO1bp4Fb3vlExt
uyS8iYIHpF1K0pDy1BsNZv1/dtOhmnOZxocglL5IeijW1xtyyHte21RvD1cVrfNXwIgtwfQ32+gU
EHgZm3oSECVewtuZnw7W029T4JJbq/GeBW3OLO4P3pqjg/UjxMSLlUeaJTWbIEr/oYDIWPe1jI5q
oPE4mKps88maeD8593pW+vYK10RFTQDj70idRyWCZk4sHVblUdRCUkCCkv1MPDuQnTU6XcT1O7v4
ttPHUISpZUOOjknauGoi16Kq5XbIYe7dlNfyQPtGVmOVukN9JmbxGl1/XXai1rWOxO8eSvkncmkK
ytGUs9EqFdOThB+k7rXip+XCKBRCeFsLuZk7QFxYP+m1bk7A15P+Jl15OJm5hsGzu4fM6FbFuC4u
Sqgk/QhKLBTcgtiWlmA1GQT3OyDndOrVw7VCmpBOY1EUq1cR/q6omBQRzahdTio2LkmsA/aoz5Qh
havAlXtKgc4WhBVeovpYpYfRTDIEXT1q+nniPHecoehK/mvN5jkNgihxYpur/c9EKiW1kdMG7li7
H4ss0OHQ0udDMfUogGxw/4O6giNJztvTM6y2aHbuZ4cf5tdaAEAsf0/tbkdYhjyZF6Iw/CayJgFT
Egxp0vkLJZvO74s0KYW4H11iHN7zmMhZkhtxKNHa+XNZuKkvBDHo/Dv2+YQvbmC6TtDiVbNpgpvq
Av3zIUmstazYjbci7bCi60fnpI6ORcIsn+NNB2km3dtONcUOchM9EJb+2Vna14UgWOhs+MvXLILC
3sWKoSxtlxJhkjAElom+wLfDGVrBt1tqak6RxWD08alo4ZV7aTvNzPSFMf8JQr7EwYJd0EJD/LnI
85qxxnlAKHFWrETFPAs2mmC6uE4Wc1B12nzw7L8inE0vgJ/fl+ysht+30SNBioplWHVhTH8ttDbd
6LvORsKmHqCZ8hh9sdrIUC+7+DE9JvxQvcET3V76drM4LMyAFI8qjnl70reFGDkTJXpzrVw4pG9O
v01nSFizjP9e2GpZOxYoULywnKSNkQDEm5bwTwZAyXgTH1UONA8stBhWfndIGL+Icidk0JhuVkVn
3+kIT+yEX3bOudE1biaD3IChAMpf2kYM4CGMD4gRjjJ/h1yNH0J9EDuYw/iciHQq2feuYRuuiFG+
/O84i7QIMTBrSihbtQa6fTNyyP9EBv93X1Gal9ceYkkSyoB0VtbTVCesBg400LpUOqSu5bPBAO1b
wMe7zswM4tzp0czVCtEpDKdN7cQP/Db5o64GzBwWEoh7xHHGyiO93yRD9MUZbJfHiLFJvraTaF90
dq4NAv32jw3gQQeazotda9idAeKwtazOPrvD4vdy5PDpe72lVyF1QPiDON6BQOmtcsgM/J3lQQIO
5SeSQTNst7KDICAhEUZOm4ko6w5RQQYGw78QK0o6nxIeQfo0VEi/FdZ/VAz3azvckTEoqLE9tpVM
JybvtY+/oybpZyThxZYORVPQ/TV4Zu9I5xZoawazgSLvcVM7ebgg9w8ApBMdJwlzvQJHTU/IRn1K
nI8NOVUpp5Al7RWI6bmmGl+VULcwfEDNPdNWFefI2rCBP1O67vsSe6hy61P/ze/U120KccJPJOO5
bp7UJDEsunDQ68py9bhRvKrm4/YLWfb9eNQ3FfpVQc4eMBwaGEMS36gemzVkO3FP5EiBumlWEQri
aDy/rQ5t2wmbVQ7DgvsBhJltdw82Rq5NMt6VH1TFm9lq8Cxnr1RgxZR4UCc3LaD14VnR9/BZqrth
z7jHYZMsngS8XnvKyInNvtaRzIUtxfMtB0KbP1s/dOHkLlsT2icVu1/qazqBmkagqzCHIcWG3lYh
/Bt5+ibyNM7L/yB/xy9IrELYQ2oFvzn8s9PtQDefZqONogBlf/c3zFrL+MLiBIK5/xRW0P4s3m8r
v826LRgNcbMcVOXdIF7Wz2pGRb79Fe2F+2l8+RJbL72EVys3zvqCCDX5TudPcUGXYP/jk1MKlvXt
J+p2FKuTu/ERrxd04/vcqpWmitVyHBqYBDHEjwN/Aj5LyX4JuRQvy3QkMi9A+AQ1bIuK3KI0Am9A
widJQmA9/uQaIaqwNp7S6ft1EuQaJH+3frzrhJQ7IaK4kK9k8kyZ0fOpCKDvmIAo9Q0b3v+dCB+D
Q4IV5SeMWJYBqgJXuZy3mZSVuM1i1uHWmP1m+idXzo2zwvjil9VnRgztVwXjHTw6d/rlkQRcvYwa
Byg9h40ntK8lg1JQm8GI3XzrIlVp1bX6LU3Fra+loJVst+6hz6Hx45G7b91XkkeuWy/bqK7XbSfL
1sYmkmIY4yUQ4YODolfKtYpVtV+ZH3Jb91bnKAFzdPnUf9A35D2ZjPEHMTt7il0Dg0pJMDg2yHZy
DbKZdI5kkGXo0kw+IWCr5SUhzhbipCkLjcsnDyjCCnmqFIFrg690R62hA0mDaHvPlzu174QO59Li
r9XarT3WY6L4cK52E85cR6a4NQt/GR5wZ/VuqYM5NOL5xMEnvRh5zxyOlieBYSVCVrR3ow/eySKk
ggsxVXDDuFJeH4XTrShtijODXgOF4h9i/t4euX7583AhVcKchBK+7Y1g41lpsggo2l9Yd+qacMWc
HuUqGSOGr2/KuaDTs6RRWebVDCfD+gXod217R3bpbnZhpwR9iY9QlrdwxG1TWOQOAmzcZ1kDUUwc
8LKXi2j3vD73kQRIv9LJ3TEYkbvv8xZ3kxp3Y6hM2bjS8Zxldcc2K363c4ubShuy0KegXfIYqltQ
a1pfdZz/rtWYzdzj3IZhlNa0oByoiGuwHWeUAhvhrw4TyZJE/2l8AFjLOFbXmPmRAH+VokZpyp+z
urmVmOAZsddKHxpbxOYwNVMfIOyaX3mKyG3qd4y01x8s7sQ0Nqeb8Kd6DWXRanytbOPAUeH0kpZn
1ItCQ4kcmQr0JIbk4YQYgMIsGc2ND92DVQcn0Cex8mwYObFffeX0WF0MA07v6rmWgRKFmPqJNXIK
va+py703d6H1l5nYJjq0vYMTb7BLsNjZ2xAeBug8b/+9pI5HX0zBm3XZsRZAloPr+nTe7VoFCkCG
ASWmn7AJf/uLq7lFm0vqrY8Dqlv92b+sbv0AqbKPBuDZ+GVbjL4yEqccxb/1I9z61VicfVOQJPBM
11EjrQSGReHngOfLiz6hV+qQUjtjKDB0CBFpCxtfjWFSpPtTCwAIa7wh29y1+HwWw6dBBG1H5fqF
NDjLLuM64ro63RvO1fAtAAFl1AC/kep97NojAMHdLAQ3aW2TzRNi7vIoxbFD+AK8WEjqBL2AmpI3
h2sayqHiWwUHXhjbV3FpRrUj888GgjDZDDSRVCOPb09FrzPvcXax6R1iQGE5b1JTPyGJjKfoqYwT
FiLzVHQlzlYlHllvwmV+VBLjNDliMY8TFsPAMVa+FXim2bSZN/odLxv6LC/OiUOsbFLEppgb5gP1
UlJAVbTbqi4/7d2YPDrJIO/y2IMupqmpUhzBRCveN6sdb3E7rikBNyQQ4OEUj4pB7vLycqh9mBDw
gsU0WBelKvoGRCs9hh68uPEn/FP4ggnW3zuYGEoe+txgQWVtx6sBYoDe6thoaymGMHk24ajl7oOD
cYO7MBwqzpa3Tw12EUTB74zFyHVPi3WZLRTzk5zBVEIYgAFBv7hTVGWp9ZvDm5aJ3JG1RTrLsHKs
tAcZusB7/DM1zvF6yxBNdAWpV+jQU0tJwJEX7YyjH6ZqBDqpjFmr9vgriUhHNLMkbgV1g27Fxpxg
vwt4tu0AZxTKrqxslmh2MnkJaM0qUpekz3yFh4sAPVjP7m8VJHSNsAVrjHwfHjACeznItAGXevNJ
RveCrfogWsDgwL7sqOCOhYHxZ+ycnbSdwHL+o1if5QlhT2y04fOZNcXj9TLDj++z9bAcFqdQpLtc
feFY1gSycod/rJCjdi0+P7cpFG/3mSd2Mg6IhYypPNJQyHpxV6YgwdGgq04yus0zZFbyp2jCSWgx
Bg7FsgGwpTA6C4U25zI/5PHhKS/652qmUXfyRvaugekt6wxgc9HPpaFJZ+BtZgdf620EjP9I3sYp
oNJ9B0y7kltOKKmM8i9gBVB/QGf1AKQdA1ngnaZF9hdtOlL0mXRcMpZQwkfkGBBu2upEs7n4MPI3
WmBX4LkSPjcHnFnLdNNcIIlVtKj9COqGKCpbM05QTAqCRMILZMSsTlGscj33SwuD7HidTzD1axNw
sWtlp51cxf/sHPFi+JgpRdScHTmHE9cKy2PaiwXG2rPnyPGLKkdcyx9yWMLCN++Mp9t2dQdk4SvJ
dtsNlOQ44pZ02QTHbhLfFiqzgzvUjq+Z2NIB4elrKlssDQlsCqQesw3vaZbdnMHaqtRhqUcmlvQm
3Tj1kutVoc8KSrQzecWLvUV1zEvwwlXXHlvBiGcchKPcT4hsdVy39F3swVa1L+3f3Lc903Ukj/Ug
1wBilT6ulm61LTsnOKfBwxuj6j/6HqBP/iDIPZLgy5WKwuiIFnV0S7pVgoBKSsBTOcN3Hde3EKOo
975zWFNaWIOTQGC7KXr0pUVJ1u8TelIKQK+z8LQFkRa/xbuauj1MeTl1xPrN2LmQn4y/fEz8fHwa
UVEzzBMkJtPKROJo+j+ASNJwVaNZuXeXgP1VPMqBDihSEZQCu8WF5fsCjVrF0I5TCh1Kg6mARaRj
tVLXbhY8lzTgHA/Jmp7q31LBWQDC5QhKYvgfupVS0gatcQJjL3735tCW+vr3pjhnqTt9GxTkkVcH
STuEsBHYx7P9QMkkBarRtB/qs8eAcRIys/swkJKDVXcZI6w42QKuu3ZqLZugVYx53H1UJdGWt+Hp
X5aX9VcW9acUHysEENjWVckJs68oCgdaXQo3AJZZtlTOOe+mH+uCdqajQlAxx75/XYzOSz9bEDZg
wQvcMPkgyxgr0om9E+w05YNu3ASRTy+mOhkmAWtUo69DiUVWWcELUW+q+Jvrg/xdQXfS5ciVkSAr
fFZOTTWzhQM3rMZBiZ3X7UfL+cFRj8w/TrUsQSbViMKgmje3Qzwk4hjdagEUapq22TogvzkYSYh7
CFHEevudvtmMigEkRQfdPe6+Bt5CqmJ70ki2Nhq/smiHMBO13ifMWFDQp9mdbQxLFZ7QDqmkHojb
AezwEseG7hI1mFL9b0bXhOvjOn2RugEJ/NaxT0wpRZgC5RxN60F7IcvzgHdlZ2ee9QbNviwFhYee
R1cUxqgvJOQcgyLgPL1vRxe/Kh/n+69nIO7E392u0ESfaEXbVUBGtphzU+Ta6v3yBmGQ8yFzMatB
6kbrby6t97vKCgnh/OMmdy2ZKDbhFhFfm3mAjWgzmuHVf12wPYq5czUUCKmH8343rlg3rUNTSROI
f/nhrVzNHPQwWo+12o+OoAjTyILDkfILJUXH+BSKYUdN7sCnwTC/B0bx3BuJrUOZg9qWsSCqQv45
koVn9ZRajbSgVql168ECtr+eCT8L2RGfIoHSEBOwI3sLLd3wNghoyiwRRTdkFuWkVVpQP1Q//Ad8
gXEUHnAWMcTADTPQgqH7Noiud65jXV05VX9BWB6wxLNa4hAiP2nSXgBKP3sc09CPu+lojlzFoGa5
ayU8SmDZetMYYguKIkhpVGnBPzy82okYLE/krKvJYmsg4XVLDaK72fjKRm71ikxbz13o9FYSwG1I
cEjSOXiUmly37FusSbblCS9YL0NzBLxzCydDC11ujXohQR5t9ZZAbjoSSGStEZTF6cN8hzkiwoEB
T7el3V3g8JXPuVgN9EmXeuC1otiQQNI34Sl/hDZnLKeLuPOGZJzkkju9PLp2Iqq3JZucShDNaiwQ
55CMqGUGrzE3yvQsvZZ9lvzBps8eSttJoJqVivqYUSm6+j6n2lOmN2IM3pO4/hxdj788TEjvuUNM
Q/Eu4wFLV+l6J19AtULBThjhc4//M74YOtRFAoOoCZZrFXcwax8gpFS5p/WLtOuWqxVgxqQf7+xL
IxU5sIKYsetg1UAeI0gqB47VaGt5pha6TPnsHHK/nxxjMzxAbW+m7hYcHJAOTItNQmNdr35kXBHy
oAzfd+1jks4/5Fx5uSgNG2iJ19/NRidHEYE606v0/eHFFuFBs2X6Lh8rxaPJmABvSoJ9ElQHdCFg
yIl0dCB4OqCri9t1879QNAlYPkPWJJnw7A01CbqffUu8HQpEjhN/iadlX/ud7fXFyyoMTs78+Y2U
wnwM8OvkkvoPvVt3GcWQNVV37YS0ZYdvmNH94HTUl90rqzax6bq7/yHEFeZtVlWhiN4qeTM0OIPw
WC+4XzmNrJPHK8dJCmx0ywryI/AcxjwcxOAkx9JA0k07aHb4HPkHrwbwC8Uz8S7GfCjVED8lqwN9
NomNoNUdEgzf4nP3gCHZRfv88HBZ3q9QsZBAab5rzyV1NuZyaO4XcYELTHmQAzd3UdQJb1+WHeaN
x5OIo+4L/8GBufF5oCfwRiQkUc/ypDa5hYGa31a0+RLcQkla/O4spOlklb44DeD9/bJq12qS85BC
v/t0AgQfL5gzmoRVp+A0104ju9dBUffPJWObXc82ZA5sK86x03dhKXuDe1DBVhb/CgHnlqFwuxqL
6gHBXHg+CHYkHVSYOrgWzUQ+Duni887+EgVuwfnDj80zRn614eL4r6zBo6RD1kANdTqOplXzSDtI
eZUnq4NO4/wyQFS+xjnkXvVlmxTxr1ROFg2zqN922PxjdRpWazOst9vmE876eLpE5GpajE7NNJdx
HZb6rIzfOKkcj/vubAVYUzez1a26NqdXdYy3gEaYeZHE/JKjTcGnEU9jEPab3ZPDmdNwHOQfNtds
OdrV23qyFGsOSl4f/83FM8dLvchn74krRlxxAgk9BCbq9Elo0wcB8/l4aD2d7/+cQ3GTi3BP79B9
HwmVv4ZwWHNL7SdAEt45rhoiJdZTBLqs6nQBI0cB00U9AK6UHHPhM24GP6EnVAi7m4FSEdJ7lW/5
E5CbLjVLKCx9Os/Qt49EytjKtX46MGIfPMNQCD490O3Rw/nIsqmasqU512S0c8XnMoSHodNRx86R
u5da+NyZPemNVFP8Zkc9mY8CxiJW6EyLipsCG30sQwcelfxFRkzqqNFQGN1jmAzqa5wkKRoa4mwX
LL5c/UAlw9BeylG/DRNF6lEK2MzYTF3kvTrYbIwpKpNDd4OJPum27XdOhB2jKjd68yZyAP9iJZYa
gimAKZdnH4Djs3ai9AMjRRrjwzI2EhDVOFnOYRA0jDvNgABv+a0q1t58XO3QI9wlIPt/YKnD5o5e
l4+IxZQ1uSI/RQUS2JIWeN+vIoHq3KwNWxeH3hkgPdqqXHNti7t146rA7DF29/08Qxv6aQEPq3Oy
AOqRGHzDz3c1b887PQ+MsisPBqCPQoCKuPKR17Lgs5WhmbVehatHe4OnCvqaYLbgCzVpBJj7nPL0
QZyMRoVE3fia4K+5uIInsdGEcRGA3Cn1IcBuscWuA3kvTGUJP5P/RDihQNeouozFrvrIrv4OQRQJ
NYOAuwhuKKSF6UJsP/ks56kXZwijB741kHtfCiTDrxHSg8ZDbuJTBm0r3Ehz9lKbZKucr9y0efNc
ch1nRMIOODQPDOiYoECxnbRwd+veeficVMljAkoLPRCgaPnhjtBPCxGFHOnl8bBUPE1Kyzp0Ur6q
vo9ketd7U+2HzCgI3fCQctYn8bzQi08AQOQ0frSQtMSd8LkdfnYY5dz2ITzZNZC6DmaviaqsbEyj
MCf9NB5dbzm8dTN21CdNlOJRoOt1LNHM2HduFmk2AHCrL1BXqO6km/fd0NU1HZCz5qIkPSoNY8Vl
xBS88WbEt2Dy/weALTXiazGfqyl73t5QmE/jBoR/XqT7GOp+udlxWSkGYftdw8lfw1uThnq7n1jN
jwpn0R5jxrWdnRlscwmkJeT8aQ34bMUbc6GJNRP9Nk4RlbfdyhPivv7mOz5oqsH3BYv4vEZuMyp4
mpgMXc2O5mR3hjnSzCYv2FewodslEMObIDMfPouTet15bTNWBnphA2ofbOX11JwupD9UGwGdA6C5
zJeuiAo10k3Xf6K0257lszxS40AXUYi2kz+k1zE68VNte567ntrx0q5sZ9lwONgjzaDt/9IuFQ2l
O7jqMN3Wg8Vs7SxQ8BEwvb4Cw5FU3awDF7Q+ebvoVGCEOowX+MCGDO1iI21a5L/6oCrEpVmtiHEQ
d+9SzZJ7sLztGokQixJ58L5m7MvFox7E2Mc5Y3jrwH+5hl50U0y0iQDgXYbLwJwNwpFRnP6pUT1m
WugNUigbknBXzjQmqOBXxxhZJbjIMrv8GABntHMp2sgYn5haadaq1v+nJIvlt4P9cRWTh+wfQOT+
/BlMe0qLZ/xruYTSaVfMgFwWjDOYZ+qdl76Pos3PFVwCFxelWKq2a6IK2k79X+fFOpZJoBSmmVBp
DTciumHd0oGvm2KtSWZ6NcruOehbml5Kx7PwoZhAlXt4gw88tE1yAO9OPaoUu0A3F/IsDoYipi1m
1IFIJLc8CfAGINNrccuiFNspdjooBCZz8+OXXvUqjbBf/Mkh0eRyxcFxs/cxxeWYI9hd/qfXwuTq
3lNbzDOpI+vEOZG5DFV2pGBzk7V/MHBAf01HBMDwwkyRVjJ/KRpPNjdtYB12VDbUs9DIVcQNWBXy
mlOchBeAR8YWarpmWFhsvIjdA79smzerAt9ti9CPtx8SCIH6ltYiGU8Xj4KJT8HirpJy6kWP1ezM
fAGHp+g6ygxVUeVmPHpDWmfwUj0Ot3KeBoHzTtCpFgaecYlDOY41BwfvfQvj18E3bGpci+0SbF5X
RlWgLbVcSSKOd+Zh4RGJIolimVbIuHaDVQ3lNWNoZg9eW5cRr0zgniJ/yX+nlfCkWFOdYimK3oqz
CtMYq3hoyQuFeCcRkvw3noCLxfDbQp/4e0JmnzMFkf389uTw3KocMFmCQMmcwo8apVLBsBs5byOH
8J3nQHiAXZYS8aZMpstgMS2m9/gnTwq0H/p3e9f3guTFSWb+G73FHw6c31ZnUSIDCfXfN+3Z1lJa
tRmRTd6cb+sd0Ygm3uDjEX9od0ikYhJuDcLSclohb3GRxLj1uINLGp2tB6WuOIW76gtFEOqu0tJ+
jUnH1s87fVsimaf+wgPm/7Okwqxucv0Pggq2Cptvjnor9XEprnNU1dHIbatBqQnjIhd3djo7DkJX
TO5BWgz/d9BKgDQcJgKRpxkBPU7kpS/D11tkx4/xocFhnD+B/YqEo9crH9akGda0v+tvU+3XuQwv
rCPUdk7jDd44InMLqdAjsKcmMPlG8MDn5LnqrIvlzX0KkDswCvVulRF4H3KBMevy+xKGuyGwl7mR
+tA3KkYxi2B7o3Rmp3gqx8jO2RlY3b2XyHUVDtvWyuJejLLmkwXuCcJ8AU0o8G3Qw2VsyUdk+CRA
azx00E2uPCOgWNQkZrypv7yui8wf/PoV6cm2BbieEVhkSqCCesrmqwREJddOZnIzZeBIGWhtNIxv
Zn2vBNeop0bAxL9G58y5ITVvLmBuLirShcp4AFQ+TVZESBxbVQrrDRv3DmdK+TOtFRnw69O9umn3
4zxtS+xiBsJM/BF6U3Tp3pq6Dkvn7e6UO2koGk9CwqmjPDwPFFobmTFRx1TLtOjIUGzsu9VMENK6
JMbAR5fErOz6dfM2JTtmhK+0LfnOa8dZgZctknoFF7LwCTZ/kGbeXyJHFjCqPazxIbw1Z0TJhJfM
U7KrmN/upXSkC9EbXHwTcdU51g1NMUiNgOvbF/Zms148k6ZMRFV3L06Bkx7c2H+WUrH4VGyoIbYJ
gBjbLhGQlINvXuqq7oV2Xx2q4EQIlJsn48GkmzXxkvrgcSAAHfeZ+OssLOA9XnCKYcefk90ZL7k6
NphEXfGkrEr+hQ3r/Q8v6rJagbVEo8YUY5CY9yyHj8S5gTzFGCN5gbsdqgy9y7tfpHJ9/1d46Wzc
a5eQy6sny8AT/ZZ13sMWTODG8a0gccZUh2SvQ7tySA0DzZcWcb6yzrZFo3lKZoWVe36CZdGRjpRw
sLih3ssJbb1hzPw2u+haIsBJe4V7ZU/2oOOEsrrRjg57Yc0fwD3MObmSj3+AEmmRh3kLxrsjCnfv
kxkfesmaKM4Q8npgXjDAat7LAmlqZKQoDv6RqmNiZBUSTnodZZbIUE1NBiCIcq9A5AswWLTPmfQX
XoD3CslkIGd9DOee+/NxAlifFSVyI4B4w+Xx8DDm030dr4+pV9Av0GYlgnYz3pq7FWxNag4kXY+M
DmlyPCyOikuoZd5zhKtmLQ7IaRLIoFbAasNwmPjXcz5bt1f1dCrWShBsYqrqyvKQW51L5vhVuuxd
mG5WOQb4hQySyrIItyg5WdYtPQIm+OqIULKcbIjJWKi4Y8/0w8nPOmBDIi8zAmklx3Pq+WRzL1cd
+VVzHgaBezEwANwOFMF2JYxqxxmzgKG2J+tl48Fqm/pkS8rxAtBN6dBrr/LdEKYaxJCAkbZNJHY4
mtQNTnmyv+FiZnLtb1scJBbBqG6T6EH554pycOcNobGQ/8zq2zpbD2+tLjJB+1ccfc5JlMVqgfmP
fl7yTqf6iXCUedJnN/X8tnjzbPGg9GeKPdWkc7y9SOt7eata1m7iYpuPVjRfWgLOR2GbtAnB/9dL
qZhe7XOwad/YQHQDy3q0ANXbq6a6hXFSm8BOMO38LsZG1gfdj5c63aECHIt84il+0zEsMyyW6Wu8
uU5+UM703lBX6EF7gJa9M5jUBcY8ycZIb+5Rybdxpt69PAEMv4oxc9gfM93wWNuLVKEdk+CkoIL/
2+G/mC0nR9sEIuUWMzxUYXVAArblP/q6H7bRQbAMBPsIGCcuyaQ6d/ZMGoDQYhIGPz6ROxDnGsBY
TLc/UuzValFJRh2wYtvDQj2uZghxqNOUtOK/udF+/77DWqtDFoM4SZXostPSJ6mNg/0DKAjsaLWl
DghcxOzOREVcv7ij4/hPLyUmqKcDtqH/ULBzqG8wDXJKZnyWopq/QtVWrILbk/HD4WEGpn5dJgQu
G/eGjMiwzl1hf6GbMm3YR0Su7D8O9oJyApwKMJjA2b0ruT5eLIg0mEVVPi0RiQF9S9yha1rwDeD+
xribLLxyayRIAoFOMHCgqs9vjW7jBh/fwAKST7qsg03ElQrOz0UxJV3N1deRTZAf3+LwMt3xebTx
krSW8asrFCyuYzNWsFKy22ohXvYYz0CPBpqrVo+Bjj0BGNCvp48QWpzJRchhVSam9ROTCM9gob14
MULxDo5mPL6S82yrkj8aSA5iSKNvGmC3Chftuap17SpCLP630AdkgAyP2xTmitU35Tw7TQniTX8m
v2E/PZ7b1sjyotdpfftGUbk7x93qFiFo+WVlq6i30Bgop+2AG/hQ+svROL0+5l1nwFUyTRGi4mb/
eyy/RGHmPkYFHKREuRg/FEBLqCEbeEy3TVdWJ13cWDASuTj2KLocBXSaRSLY0fl/Er3eebPSsHlM
48o8It7R/PlfsfnrdAhy6AEfiF60RgTBEshfhF4JgmDXkG0mBRwlBVAQaB4Q5azRGId0VABOty2Q
7duepHlDOBfa2w182hXRKwuyfWCkeNI9dpybNIPpK1qDv11mq6WckH1jnQlvICgKQfSEyfYyt08e
R1XgHYd8YwYS06POjzEWBDvzvFCCTN4E5n/6RCyGAmVBZdPiH6+B82yzPBHAfJmv6n3EqiqtZDDY
cMNlGeCcYxVUGJ9F9dx4IWbYWLLjlXD0CWAeJ8IDxdTxwIxDL+wEUOclvqmDQUPGqmKCpkdmdP6Q
9UHeXouOKzaLoxzhNUoq8PypQpA+Ey9uDzdokzi4QK7UsIimTqhKhjzZ6g41lxfYUHQqKxEntJYb
gxNhLZAeGnDDBd9v7IZZxSoT4REQ8HpMSPgOVci47HV793o6QxdiBUsffzE1y4rB7yutdWaOQf6f
sFT9OwFg4CoCc/IvS+7DydSEVeyTuF2cuX6jXoRfXMY5IFMkYFpLLMPmhR7pg6AutD4A/9bQ3Pbt
YhrBwfyipx3p77spd8u4l3qxmZZsUN+4B/zRZnhu0ygaQjLmGFTocSGE0jFpyLg6RCeoTeyhvrN+
jH+fPaSIvq4Dmakaw3HVBWy4eFFvW9E3KGm1AL2tZunfiaSYxbUrcOdQO6JYyX34q0QMgqM7WiBT
e2j36VpKxGyxIJPwMvMAqWD5xxjVfm7/2OB3nrH2EcDfLtuFVYViLCjoJ7zNWixXx1P1WVQ4/mwv
XFgqsEDVsLuUfXXW1l4JvqphFpL21DitUjap8D4eIinV5qjUamvNGWoL1+MSSFnzhS4pyR1R27uQ
kngt2pELlpxxTDPNvmh2f9lNzfISpNp2a7ZQMsrFxtzFSbzZbqD4osVSKPQmHoxZVRgMDRxk5fWx
mX4iZGyKFUQv8PMtRvy+Q9T7S+Bzy4Nz/JIeGkNe1uuT8u9TGqnUJISjAwjK2lNi7+x7QGGyjHSj
cZN3BTM7zxgoxjKiUULRsIRqfSYwT6qg3uZ3v9aRZtJL/ez7vcQyjR1qjMU4sem2EORK7rCfOSt/
55eRqnVHHOHZWYc5cxzWZA36lYGrn8rd/2Mgxpu/kh6ZNImneKDX+Rqm4XROa6EJnMv89Cgpbju4
XIS0x6F6qO5OLAKHN4FpA4FaBk9fz0BelZGAgy4jD3tBxy+1DrKYb2KCsWVZDwLKJnKiKR2xax/i
/PuTwZdnKHYmVALwciGlp0XAih6aySRF6JaAsWAWGgVXdWVwQ/DXHvspTWA5jKAxBzfnpNsa7yPC
0z4HU/Nt7zRxrVeiKl3qKCtkhNdY0UfOw97QmcPSai6t06FJjese8wIw6AjFm4l3GbEmsfI4Jiug
+koWopioQCtz56yMmasX31y70zzr27O1fSAhGr7QoD9o1my0ymk7CRcMq3fBaONyBtVXM3tO2JR5
yzV+Xmnh3Q6iG/Z/kfs92NQdYp87Ny76LNC7i6nbpJaG7654YeS8771Y6D8mXByvbBoqPM1PVNgJ
8EtUJyVSKaTWL6BGepr7qq5IRE0hgi9SOwnLpxrMBy/kLsJojO23kIxSytheqMd8QK1h+0c+IIc7
jZr9x/e6A7uFAHQ9IDT+n5NlAOIYm3jXMaS16mfMHd3gvYdvWSkfj/W1xKkbmvubfwdoZYby+70t
PnLpNlSi7xXPb4q04FakWcMcGeVakFJovdrSum9z9ZMMoWg+rI3jTLaXE0hu3pedGVdP5vAcmoy0
8w35uIZq1Usn7YkhK/odBaYc5CjC+B2sD8/uD5nk0CfT5LlqqdfEY6cOiUkhv1vfGxitx91vE4pb
00k2pw3x/iqiM74yrs4ZvCpesKoByYTsG/oM1UFhDgb3euUpPvhyWsZZF+lKcDTltv0RWakrkNVq
POaS2yYfRHCdw7jfuvKQTNcaBiwvc/MnE5ZdL2XV1raJ/4MCedzT6tFrXzFXHJjP474UlgdZ/Jta
mOSkrCcSpzsMYqzc5QIrdRiIB6FYOC4yp4JtiELjHBtXJlDc8D63d2Db9jDHahgX8nFMtf0Unqiy
eXmdJfq75IyxzI2paB5ZtqwpM78xSE+omwqujyVrD4JoiHy91vpP1JcP3Fh5F5AtsT8MP01xvcex
kH5FSsyccuPnluYH7RAJK5GKe43ZQHD+tg+xDzKlLJnfz/1f4ZwOjP+5Vc95PS0bWaHHu3UdDoIk
87kzQ+Y6J9JoRGT5261p9K/iZOuKsm3B8b7Bn9lKPxGdpL32J9aZffcUxmbDKdpEFmQyFfFw9eWJ
M/wTQPiwba4isqNaNZUYWFLHIWnjVQbACUgGxqesOgp6C8mFbz7RptPvmg2ajYAfCkDow/1Ym9sE
JS+h81H+NUl1CL/H6BiqmjhhJ0+h/T56vbm4cFnIZWjvS3JssrnRSaBJRbzb0LuWV9pa3qmQK7lN
xI99fRZnU0Lnxp3fFaObW4/kANZe56f/E9rmeBQ/iGk8oKcMT6gxN3WexO9AYDjnXd65XDq/gDuL
oHTabUR25+mMBRon+lWsDjK5MI6PXqACfavv/eCHSWyennrajstxFIMAowJi3FOMYbZSrRZZnKYR
C4Ti4EAiLU8ulMNfNFaIgj/brRs/0ibxZfoaoF1TO/whyVwUN/v2+SpUttAQzuwePQUgYB3O+L/D
FlgrTdFe9B1/T1/Xk5kQ7ypsT7Uum1U2IP1bPgtUTTDdgZIlStmxwdCoHWh6s0l0SH1YVSv5OOT4
/eVGGo52+kq8jffUM1kbmxB7hjqU8+pCuuvsk9F/zbh0EkZTSPujKL6LumbQgwAashoRmb8LE3OJ
YhKT3P2M4JAcLHPQdJR91ENBah90C8SBNgeIiUxESCui1FUxa4Y09fkMe7XWfEq/bKhP7LEAiMe+
6icsca9+ngTcmROc8M9wyiSEghnuQpaNJIgSa1LTYzNu1KtH1wsA6wE8/hgWdi7EF1IlFbh1+dhq
rFpLPl088oDGh7sQDNxNLq1IIgKikItRHpg0DuN+rl0Uec8DDfYezfnbeAQbuL1WqxPrYtxpYlui
g850AqMogZLawh0TYS4V6Nx6D5hUieNUu5WNI6MAvJr6QWrn32i9SCfk6oDgcrcqJ8EbLGlnfQ0j
Kub5gJiGHs6REBJ17TFWmmGu1QsK43ldIx7IkKjMQJNDHsfBiSxuSxf1K4zmeu9M5AWEJ0KcUfEk
uOmwy/iMviiHuAC+Nm3cYt2Ax+fcWnyPRlgL/ldZgogBXk1gEtMI3VPTc9Mgn2KQAYuYzgp67qUz
hoJjDnm1e7IJqZyA5lmUMqFReC9+CM1kZ/bGbYOVNAEodY/SJ6P1Qbl3rMHpRzCXOFhRM+JZlSll
VprGVIz8GlxBwja1rTuoOt+KdLe3xKk/snd/6++XwUi2sLMn3IW+9LkTgfpzI/MkR39L4bYLtcEf
FWC70beImYBdmQRrzQfOJlKr65MB+Iofy0p0ivRFswXy6xwsGfJm/S6t1gjVsxrEVMnz/NIN+FFb
CgtSZJziUOj1TeHrVdYSoNFRCio/IQXIcQIzg0BeTHI+U+NzmUE4p4Chiw1vop4QhsjwsdekPYAB
s8k92QlrTbkWYj0hiNp+G56B8fyM14BOPJPH/+wFFfft9ePHecdaTUDtZttaM58H0FSum/ySI99c
Izt2eLtA+BCb4xNmr6djOw4y9OTBIG4nwBaX49Cbe2q40zdbUl/PJW9tsgUOu6gfbsFA4ypn4kz7
bbLMUqpYtgmd8yieSPW+AJFXD+eS5yTvd+JPRttuOPWmupKFgtBbwUqzrkpAheX8TthXEOD7QbWX
YYzUUOadlubBA7YyCxkGm/lJhvxfptqYf38g6tdmAU1HUq6ashK/rj3z57XdgsNxXYvD3vZUckKC
rWxABI7+d3bfVHXMYRfamn3TF8Q2AYVGjf9IPgnF+AAzBXlJjXcC/Y2v0tNlwj2GH7rDU/66lGdA
DC4jnGRHzV1+SQI+Cbw1mN6jAyvG1QdXIAcr9OdMQgjjtyLx0E0E/sC41FHp4CZw8OwBj1ZTDLnr
19d+cI00xmUwyFZxpIc+619L6h8Hih47TotNOfbJ+4wwIYBZQ9hpi8wci238bjdLFtV9NhHq4AGQ
CJe95z8zC90cEg1x16yVD06v8VYDdOI+yBArwH1UwM3jAPLuI8OwjU0Y3mYYZN35PxND/VosBesI
odOeX7XLB0/pomAG+2ymc8ctbcUHbxj2dGzUg83tql/j2bNtNvmNqRTXfw+c/fDaD6t3VDwwys19
r5l+uyZycWO6OoOumaahQ8fZSV5JanawCWrlzUw1frHd8l2OmE0dAQTZpJn7aO2OXx4WWbWKic63
abrwSw9sNzZghGl/2s0MchaihxoBRITi/zkMD8sg4YluTDWUfIjO/WlF4Vp8sRu+vXVe9W+d7zc7
SNe0zKrLSEAwpMEXek4fG/mM6tUAGa9Nw8s1f+ktUB/iZo2SkOhgXM/ZnummaLX6iQGSWfTVejhO
OVMuMidM35daP+GJoTviRrWc4S3zW7Bl7rXzikJFTzPv96ku2lJ9Aqs74Hos2l0eNDSMZCWssyWo
XMFJ2fX1DCJhMeQbcDoo/BBrwkDfAkhUjKDzyD8ml8xCfyJVzQ9HXubccE/TB2CSrDclJ6ASJz2B
yx2nr9hXqGUSVgweMOZnAzp8p/890EehdjShhexjvVp0TqNi6ZAtjNj8gDnDOWF+AbmrsJNe/+/1
XZjy1xhw8jwOhG35pwkM4gQwWnownkUDkUIoj6FNJUbDfr+Key1R68KL7i5HaNlzGF+XJJa9cFp9
y3klo3O5XKdfvdKdAMgaIPBdXAajBFgg5n2X+oMFoA0w7WP/yLQ9V5T4ufPf544pYtKOm13LhC/P
wIqvHfZh9znypmc+cK9CKyjCOYzOBaKSZl+cvklQyXGipjR3HSq2XkJKyznFHY2WYsRVXLnj2HDE
tXLzbIXLQUDR7UNm04tpbNa5GB8voK6G1m9nap+r4tyoNTREPg6FXWU0mEm/z0xyJbhZ2Q6eisZB
/YjJE4SHACLIQOoyNfQZS7K9kIlCxkGdEM6ANedSwcSrFcZx1q7i5srbt70tuQbut0GPX/yAUVBK
LM0263gXmqTQ0uCnCoMuYH1gOFwiwrhC4amgB7QaTrobJLb1iD+fbPWHkxx+HHF/1VPKn8buewRD
wF9z+pSmhEewLXPTV4fNlta25j/VFMESP9Wy6IqM9MEOsIb0qxfCD36QA61xwoaGoqbV92TctWE2
FzCGw0nJ7ecCX5Vu+IUDYBNBR/BfWxlX2ad8jXuScyw5+K3PxFEMA3Lt6o6I+4Bt5czGTgGdDQCZ
+FEe96xvG7wG0WH6c/2hihv9Jey0e8c8EkoszcZR3UXWhrhlhdPr1GM8iCX779iKHLELcrxeE6X9
y7EJ4mWSzf0Cx8QkCVXF2rsokYDX4/9xEvTot7XzfBNFJLsvpkZiti47gcuPPGjr47NjvY9b/mVg
lp53FV4oCozwL8BwINDoCgwheVCfhqI13Jlr8jsPuJekiZBdrpSawDyRo3vs2bsQYFhys8o2nNPe
kKZ/nWfBujrXIWmr4E88IDkEko+xqf/X1NTRwSwoI/6jfgbYVYyOUIVZmMmnDwa0wIuFWEQTYqB1
NhEV/YU0bwU+0tZfY4hGTCdSbb16lv+ImguuWSc6Z4n8FaXUqnbFCWiq3GmTHfR9l84pBdX+rPb+
ciqG6suoW55usmb5eGAM8ALgR81XBpOqdNGuMI12WJDNuuTUQ1Po/v9NWgg3bvp7xxB1z4zz9fHb
vkp3LkLDENOBbesgxPa90atZdJxziHz8gVEKVJmhasUQdVuQ966pLMex6y3w+uTAQFELYLL6cuFA
JoVXbYnGOcMwj0T62eWi//NjhPzOS5wuQ/rFeLhKot2oDDtA5VjKiNXFPjWCyLJRlmo8CAO+cDr7
keDtI27vAcuR17FJU6SHFS4O7LdocwufzKrxLtvYsdGCosC18Dr1fpz3ge9Zg4nAyD3Z0ME/sL0Y
VJP1iuGjVRLIgzRHEDS5F+5ILeObwixbKzummeNOZhvyHi1zwDdnkCqN5br/yrRKIuDEIhS13tob
nJ9wYbNbVzcCuxzuWt8Gn44FNFAabnPXFbD5Lkejyz3bmbXClTsDR1E/5LmB+lNRS1EZ99/3WQI0
6BUprnG4ajprdtQprIktYQhNju6vniqkFTyFjdK63+8LGY2ahyPNLZceE02WBG7wth3Z0FCMK0fl
uX8QaKJa3GlHEuL9i/Kc2doDWCwDe1UpFGYJM5K8uu0jT9lRu/V0tkwd0T/PaXuxjOfoLi2ESnXC
yaKTW14k7+KZt4enGpKSQ8//UgKGtTuM0NnxzL9Ids4xbHP6Uq5v2JuDq+kuRr3RvvtU6eIdR+9h
fwfDZhGmn1A6Dh0McgDSChIkxJgB2QypMSo6HCZSBw28JjRsnnNIu/pRu7axPAee161lOOfpVA8B
f/aP01u6Ldwld26qqSoJ0pcC9/u43CwF/EEe6W7Sh3SMixGzD5a6KAeOoOCvicrB1Fut/GZ7lnyr
H0Ky1oFZBmB4shHz37F9vq2TyJXGqufqhJbmNruhYJDDgyrVqngAYJ8CmY/0/z0P4oJW0VieFDT1
bIJCXEz/qgyXyMTKaq7W9anV2gq0naNvy7217XedSvTCa6r+2pf7Nlml7t0P15+JWD7Azppa1mxB
3gBYOHmzSQOupppWaovBkrSF7go/8qeGaUkNkBlsVwJQns+wxV2FSMqXL9GeiAPzOQd+nhydlobl
6SdFqbH0JFRF0vDs7IgjP7BvhIp07c4e1DnMCiIEJTVDVKfhz9/tTRkUBEuIc0TV4LssIg0oTMFf
HEccbw5G9IMbzcPvF36sN4Dv4G1CE0Lp67/Fnuc1q1OTdeeynttWGb/xvd+KcvfvWFu3zhGvZ3nY
g8FCWnHLYqgLhPxRQzwhB/HWEggsuJRmBBnX46IA9HbOJnjcA4ci2s58o7HW7951tY5/kif2kMFV
8emuCheZx4hOUPU1KiJ6VD6Ib6YUbWRHf4oH0QeRb3aBLJ3DO49VyGOqjrM7LB41HqBi20l9wBtu
o031O2VFP+how5FOvzcQm/H/9WJuQe08Fa/SYv4UZcYFdIxvtGD2l1qyjPkDgzB5GMcERqMwfKxf
lzbTU1Jh7z58nfccjME+TcloIBpr6k6hMFtwGMf+c/6yY4rzC5sy1Em/DP9MxNYcJimatOvcNNHn
sYjZ5OWGaBlazBjVHZtspiCP8hn9X0mZIFs24GsY5UcfQm3eZgwA1bVi/jEXttza9bFNTo/Pbdve
HnH2ZHWe+amyMlbJeUBJ/pab0TPIQtDVVxMeQZ4BOHvWqvP9uaYH4FOKaw2IvFr+g7usGZD1X2M2
HxA7yvPS1LqrLc3nV+IEb+eu6gLZfqUCZUCEfQCNUrXQRxNVBjip5jybLnJ6CKHdQ+GMnmABvBdy
KcCewN4n4xZQoVwIfT28IwO2R0hgT3fMQTWCe8FTNW0QuckWW7zQunJEf3V6rwclYyfjVG2XhUzp
XKNhlrCHrp2L85csnz9X7+YQHk6TNMyGtW1HhXgQNvNogYPcLTiMnxO3XC/BqAXpIzREq8sTmsXG
COqQWtPkYlHU2nIIPEpTSljQL3yDu4jNezk/VWEjMN0P9Q+iE7JKMyHqfbz292Q2ptA75kX4ZAWo
6Cf+5TS0JvkuUK1LEAljwIAQlJ455nF7I/TaJxRRUnvaFmZT4igVv0Mjd3IiBLxun2dhYiVfe0Ok
iIpHfYAuBoE5ozxTRWL30+R74p+HxELImmZ9JI6bQgN9hQadhTJ4qJjHuHJL+U3vfB2JUA2sx0DI
16m8lKQys97zZuHWEZBx2lfScpvkTY4CSCf3WCbkr9TxWLPWYGF08CK4yG3q9NFlOq8rsR2MkFkG
b6kTXmhvqeQXTC6EfRLIhwqYYRhMoGCj7ExASqYr4tsbozHDu+5BRn2bbcLBdwmppHN2/WoDFwV2
5wBNtbTtvYa2ZruDZAqNh1Ar27AUhG3vqQlzu3GHUltJDwcpD2aWF2ytj6uL4z8e9QZkvbuZWow9
gPBuJ7wkr47cxOsUxNqlbKdxw3hl6JYwZJRdZJrs9sFfeDexqcWXRZJ+cgYCT49lTrhnPHAM/3A7
8bb+hkIBHsCeQgLzKwtWpLZt/NJ3vhW8e0+1gczmFsgx2cyT+XIgqO1WDFrbyaqXqNJ4omsRYnML
XANjr7Bwmt9gdYMuHVh3FthBG3dXHmIETkabFAp143T27w347e7XM7tueEHW7CtXMJb0BfCgLkcz
j3LQ4R2+2SKL3w1+CPyBtta4xQ7oHOD6bpOcQU/VDBpHIiOvFtUqBCsnSFS6ZAAHBxZMvyu81Qnf
f6EgDoqab6/zv8FEca1/tjFpgRGZCxIwNK9N3mu6tFnfNeQqqA6HqfUvljfoAckd0XThlnT4sAGL
jJhd58pCuk5Y8lTQF73/rrB0hxOO4Nkxj0KjG9IN8xk+cG7vXx2dKYpSOEvLETsA97hIHIdzk7GZ
ttiXKueziKAFyOX0XLhRfhGjj5WjA1e1PVonDuEVaZ54Yjr5K1eg0uAavI1sr507/ZKtp2yz0pl7
LtTw/TPk2cNGNV7W3GeAMxtrFQm2Q65AsUMH6ncu/PjHMbIfIqBB2prCKlA/YucK7c9XSmWo2syW
gne3wnLBOR4VY0dTCGBoWSbW9R+eyd4c3yr6eEb/QSsiD8JxRMMl8ab7GosrjeInWLm/d4rQKM4H
emkJdw17NKvMdlGi/qCdMJYRfeaXwf725Q0l6nG6jYiE7szIXkGQ1ekFV9KZEGXTwCuyrTfDyXJl
35iVdkl2axUmHwssrCU+MMYuJ873tCnQQTjv6jaEIqOvppDxnrj4P6l25WKDTmdswZ/KyzYTqltT
7nphybw70XEL8OuGKFGtzben5sMX4nxL98aZ38lsJygr2Zn758lXQw7toYKxCjOylc1nVrKIMrB/
ojJqgYU6euV6svbGRTj9gJO9aRuL1RVX4qSpMLsgxHwv8EySXCHs92J5ir1CSv9vkGvmFx6xvqyn
qdo5+8JfT06Ut75nZVYynkD1iimqXSxcOgBIEjELnZ9y1R9+zBkJB65hcbPMjWdNP0SJiq5/iVpB
mU0A+9EQaYAbti4baWLCUO99u4kkoSkTcGNd0Z+kqdrLw03KydHXgS4v7TFK4OWq4v5Pt9bYHWMF
Qmr2ZRBIvOi6arVg3KMQ9ijz8pVmr0xiHOgzFBXnQWW58HGf/wZ0OinlfMkCNEse9KxBhuC+x6kA
U4i9G1mgE9zx8oTt83jefBKeWXjwNRWVTkBnl+2WSKw/ZabIHQj91gWQM+KqHMhRsD4GHLTQEz0l
WDM6ZQmgy1bKWgWKEK8GkJpnLoLeKdnMkUSE3fxsgPX80Y4tgcLOm5K2Si422ltbQ9MR/sw166rJ
jccIpOITUs1SZGjrga2eYTNx9UmP4kjHeS1ud2uIjg7OU8cnN+iokHJLRa+YGrdxrQUdYSmNG6YW
t+xssxVUj8KH+u5qqImYh7gUnpd4WSmhw+np6OEvogmSZugQEyF4gzLhwwHTIUDIedrKkYiSkcHw
0ht48+qmFn6Mn5sYnKfBJcvavl70rQcEYSNO9pAA4kK/5ZP4NvIWvlCt/cNeWz3k1NokMstUFe9v
OVWncF+K76mytBihflfKwqim8EHLbZZ5fhcb/1qOEG7JTWFrtzDYzlio41o0Ca0OKO0xtylQvWly
oR9wTNvJpQaHFk/do6wRz56aaMV/Q5oZYqQZuv8YvJiVKzU3Hh3NWBgMPSl5YFzQAugZiC5Ynnlo
gPEUyVE7oooD7mCCWtyed26XnG2u1K2EgiTXvd6SGIa8395z7ivQ8CIGR0iDe8Gj0qEK3wtsEZGK
goYexuHZU4lJAv4aoxkbtfJ5HWqw2q/6c9v9nCYNbNQhagNAmY9FovuCy0qdzYsGTXSHQWe2WIDa
isYx/DPric8HMBtWNge4xCGvSswqCSSW4+rBpg4nNaWGUtRrebOUvTxUy2JXwy3qt8Hl0UDGS7b5
8Fzb9N97jpJDo4rG5QIEsvOiXmauf+9abL0iqqNeWUQs7Hn1AxgrRhew/MeZjdbtoQX4CxYM0FFg
DYxNevBUxRLav8PNhGSGvJFRU+AurGGf0DakmdKzcQvYHf709rUDUyH5qofP+Vw0rf0NsD9Aozq+
bvRoG+CBCXByPAnIGBR8ah0miVvSvJwAPzihqt3wBcYS8KLDWVqf9G/Ulpl9+9FFfPaZMjBA512/
98gnXl5lmSQfQLuvMqvKPWEdtNchwaE4Jj8kzSRRlJfLUN47PWfVWdmH0TgbQAJ+b/+R0ejtk8Ev
3fGeaJGIJOnRMrG9IZ3VkFIDTyP7kWWck6dyd5lDOkti9X/5TCeJ+ryyVeP4++ElT3x5f4TeOpFB
uhGXSz1Np22QzZxwTmZM6i6l6vYvLnviZwWWLQv4DjLUpHBW1HiU/TX3tkxOxYxjX2A0Z+G6s873
cdl3GYb1P4LS6ITofuueDCJYsxaYjUJPSeAOdek8fdxgOzgcbQnmalwLPoAb6K/wUjfzcqMQiP1u
TZfyMSL/nfKhuYUE/npq+LKy9qDBrWM+BZ5ME+w6eddiShleMDyrvJeu2+rW8na5cSnyOM++s7fJ
LbIH2M3L/7Roo8++KUfyCguSHxxscmMYb+QzTc27OMk6LmzpfOkgInGVGlZ+nFuajGDKu+h0ss2Q
0KZaCsVjq2HWp2zgBqHUCI/TCfcGadkBybIlKdfWs6gkFNelPWeF5qGLhpJI3+uZLc8Z4r7UdFMk
n2uFImhzzlIEDxs0rEW5LTPb2eqdiFJb7iCtCpG990jCu9qmOhlqgzQIVeQxt10dhL4Ph/DBhzI2
LgGG3riEwSn/YC9koJzUqukPyBd2dWMf/0JA086UNODNYPKuReFB4iCzeyCyk4RjWgwbO90tqr5Q
jxTsP++0J1uJuzjbOT1pKFc9kQ7bFhOZ4tyUVDsbc1DFSajqvjSNnUb4m2RtKVjE13lLR7FGlMkM
lVyD+MK+QQs8twmyZCMCn5o828aiyF5Nhpd+tqZXUZvX3kByUk4BstceVX1emlsEWN8oIzp6cKFB
mhDyRrQrIfV9/D5FZEPKMrRLc+ePOtPx4zel/dYMB7c27fNs+dgACg72NCURVaS9EQ+wTDa1AXwK
39t3tyBCn5R4qYpU8/ZIi/owV0pOO03GNraKTZfjzF4pAMHuZ2KyGAreA7cEbqC1svA/RmwO1sZj
zz9XKmrGN1B6fvKfe/S8toJZvhkidQmAbamPxxKbVSaxiZKq8M17o7OJJKVF4/B9NLnnhlz23lwW
Gp6056wbAmeqpnZSC5TiWmgRrLy1QXljnvJXPgjC/H7tvLIkhTXqmW/YkQ/zRubYrlF47dQQjemk
sVUIqMkiDcOwFqzPPOTn7YueqefXXOSpQftztWLLgCAkzjzSaq2P+T18Vj7SEQ+V5mg9G7MFQR2l
1QMzVlP7Vz0U5yxDkEUuFkeDUVr9lylA2WujdgPFD1MqrlRdM5Cqhk+gVg6jigfj/S7kNqnujy1I
YJJr/qYOh/2wbpDwELnoDpgkbSdyifZegDHLQH6tna7JucXZDQo0+MFKK/fHbaTIEcL0VsXg7BF9
V2HP70QhxO6SErVLvK2crUXUK1T5hLi8msPOsWLlW/usaX1FGicWcG7qdRkKfHiXyj2hgeykmbbJ
+lytU1U+++m3hrRXNgQ41ztpY3+VR1rTlKfdIUxCvBLLX/c1Ct2ZX4szAE7A2gN7iu73v7FKsy3L
S7q+2xI/l8UKvYakv5dIAGBXPWITN8l43zTXdTZIUUBkW+Bi82F1C5lusP+uEg4NmNYSjtIwguF8
UCBtPGDHNoBzGHBUg1KFOxmBov1gyhgNtbOhiL3XTanxGzzEwDGVbube294uSmjauiMF8rftLCCD
qxQOfSpR8jP9sqHsSj5bwsBSXqy0W6G6vvTOq70XEtUVJ1G9tU/tUShpPKs8SWN8QBaOLmpVH9bU
4i8AW5F030WH0v/VI3hd3W5p5l7m88uNJuMZyUzdJk+9dzDOjVrHRXPtoe/kIfk6W/KzpizLT+ao
5l7wSPpoOc2sYqP5DkU4PhwgqbzHG8bu/kxBSMxnaSHdjQlYXslVnvxPxSnl1u+WkSgkI2I2LzAA
kmglCH7iA5v2t1+KYyzVe3dcmsLseV8DHSWKtS15I/1mTAnKQzILPngRQfjFNTujh06YkD4fHvmi
UZVeJymh23r/sSNvwW3jqhejxdzT2/uNQ7OON1rJhMvK+W+0l+45bKiRz8b1ouMbLNuByyNnGB1k
nGbmYQozZ5zbWXZpOq36cKOPbaZvOFyB0/spaiemutNPg8xZgKr34xMvBEc+Bo69hVQZFXJb88p2
d0GwPL9zZRa4xx5r5XSvabzol1Lo42QJVa6yZvm+phlXeK15pAbkMJSGo0wcn8irm1lMunT8RK/g
POUJs7+7QFm1ybZX/Oqqg9AqQie/AyqbHFVJy5SbLKYw0pZUqJEwjqFN78exkfZHJi6UyFaCXNPb
7D35WsXpjanKE8BRJq8uj8Iwi5/nD5Ct79r5+lp6YjAkHe8+bNLyT4JPZFOZGCCIGEENJOB1HtlR
ymsbhUYEtYchhj0QhdIxhBBpgeHZ2t2WkADwJXDmY3w6pd6v4FwyJaoVbDRR35vN3/bKLbna9/V8
gRKgyKl2p16+V7vNayhKAh4KJjrECoHHpuz+nmbd1hjOn+Oky9KWYf57Nx1JXuk+58VELrKZ98ye
GRX+Cf8urF+lfpPIrT7/JfVWkgOnFhpJrv4wJ97GyMZy3S6PQlMsNvb0TofyYbB5uzrtcLZUQeyV
IJH7rNwjw9YfnEk2nCt/5PsCuwaGP32Phe0l+SqNWiK04k+Tk6LFVBNf9C4sg5qrwmGfk3qgNFQv
Ba7oUpz/HPxPpz/Nm3PQDdCzLashWiA1afeuW4sziKqberkrR65xz6D3qN0sYlIzqrc8es6651in
ADtomr5hWLfsve+jgmcPS6osaysbls1hjLcxErZN1JZzeIREAcd8kST20WUzSFzPmIjME06XJe9H
CYcsXUj8m3ZduUgdzSfY/ZyFNpAgUxoCke4XdCrucLIMzIJOk6mDiBIE9fMcX3bTjeNqUNliw4lt
tjbn+UVFCEtyAH2UDhsPWEeK3ht81OXIMgRLJRIY86JbijEsqhwGEPhxq5D2kPEDW3G3uJF86Yf+
IwmA/QrGC/oJiDD9dgcO8K9QzJr1W+UGPHUVtsIPBWcaGe0CU+Eay4EXsqhXUL3Xh4+t6nBBHzRb
pBi8dWjk1bt1NtlYzGfwvXb/sbqIDgVCusVfgFyvKkvt/wTOgZ+18jRWLrghZIDAdu7UgfgMYGN4
3SXoIzn/MOw9RDyLNRgWAmsuJTBAl2oBhepxfQE6JZ9EpVwuEyKuD4g0Ap5ovAaw0xEvsyZKeJ7F
pGwJ+UHCguIBGtSmTeGYGzulkAfzLCcDzVHejDLe5CMAcYHpOLAOdt6pDnSdexxtiDsqc7/2XNig
BfgvAhuycCK1d+iHjsaOWaJbjDxyeGsG6FB9r/X6crPPSsN75y6jgo8Ee44daNnnXxqjl75QDOAC
hPt/rDGy4F9gsNRJC7EMAzcWa9SYyaGLbretF/Qtfjv8bbwErrSoKBTWdLa7RMv8k2VZJ/0kt1vR
/0J0nmMMxyIS92q0dNbCgMjr6jlo5FaHi7HIY6fiAh05cvvmRf3OAVNi3+5X02DUuMLqoutXhjGT
kSbfMcurWwVG0BJMbSruF2+6tExPl+zm3+1JMaqtw6ewZWDzGJ1eG9hoW4t6t6MhyPapud+NTDqm
+kaFyO4Sgfdxr+dlQXOK1c7NexGbvUBAWtDZ6Ob3aoiT6v/KzcHy8fNgyKKQArCDyKTojwbfUidt
7L7/Vp3iNgwSGxnZ1KYSKHXwotZP23Uqy3j+BhXRAPGGtjMNBOkidn6OAObuhwWxz0v15k8/54s0
FgiPaCSkj5FOUgQXINi9bIhHdeoMMO3nX4ZrB+1IQmp6BsuZc2qPdU1dZF5YhN2oWitxY3WSZ172
Jpwgzwfzols5XsC45AiZz2e7CFB+IdGCQKTY0uQL6RYDr/82rdJHLu3aJAon9QMEHz3ngDfsaR3J
Pbb4b5XxCB0bNLDO9ohkf+gt6AEuKeCagBUeYeXFZa8VIi0v8FNyZ3UaxFSMPoMrfpdGSzWWaDoA
FNWI3X1k927NrakuhQLKT41Gtc+MRmyZe2LTlQXWpaSrU1uJaNBwPjBG+DYGn2GKNpaW1Rw3t7qc
4knMBkPu1dio60aRb1eiGQN0ML2GNRvaNJEmFBnNs0IICZ1oRCDwLmKbnI71JxDGwCTs0jGloy+/
IC6i1pOdQKuqMZlzC+77WKf5d3BCVVedBwsud5RgXNxtVnKckLR4FaciXAOQWaJctuITgYvZ2nD8
z59WYsuCFgpw0i7gJKn029hr29HoOcgxsvUfqclmRbz6ZMbA4VeRaI08HB6+Pr6SOERopWWRgCvb
F6fuZ++5+h5wwq1H50DdhLcS1Z3XI3faZTXiTLBWdRLiMW3Ge9nPVM3Gn/h58ASAG43dtYohzA/Z
pXG+DCUUMRfj+ljMIwgAZK5/aNAOR6g+Ol3I803szDuK/ZgFrXf71z3NEtFRKgD9CT7gsX1hNlKv
B/6OjAD0dmv+Eh6+KG30KpYjIJKkDHeZTYWakkZdHIWkkymHjUeFxO2pkypuritidLE26AUuBmOR
Jb3ivENbTvNcDX8shdMfslT63AqDJv4QyGAukfLym2qNGDyqFAsunJXugwdWWI3wwiC1UeQpCZwV
mQ0DBrLxVTo+MYCRI0xa1RM67AQqsgldGVMpoaqOCTlfsbSqFJFWFiLNjInDGRsX2i3yfsOQYmL1
miVNz0IOAGUx28CmpVd/UpvSJikompnNLdtuuyHesYmCiHwoN2MlpAXBKEHByLvUuizDLHVcsjKI
p35fVF2cVJ4GuUeWX7RQbLL9om04520+gUqCKPNtkJ1qvIbWYKRuNPM7NRTyMS/K93WHv4tHLfH3
BoO3bPDpaHaFWxMQRzQh5RvSu2mAB7F9V8nmxWVJIhVcm6JXm9C3Lyuz+pXWEBNzx22Le6aJcqZR
cFHaiO0m+jfjf9yyKb/u0VbL9aDzSJzAH50Vuc00VAswPcLzOY1GQQ5dx57k8VBOlmOtrylgU8uy
ooRa8K2nlf31H5XkQmUqQoli84tVktijJBbf7SWVkupqyOLOYhPnIWyrrlgEPTeQgZW3BwulwB/p
vuja9SnunSsdbmrxg22isyOTOo73uZJ+biRdKvyH/R7GI8iFxRtYgDyrcz19+vswadEsDW+aqoWh
La67U4z3Ll4E0lYVkQk8DzpexSEXKgOKG1BXvOhtaco3SZXQ+d60IFolSYCAqsrScvTeXRzsxwR1
/aAH4g7hbKtcKXM7vOSLvp4ItKTmS0QdoYedju0V/0XUDSqCrH0WXfNqUs6xbVRJN7oQvdFzuaJQ
mFRAvKPPG5NX3uWmuAYCPbu1dZolKR82GSWba+/VmEU0BCPPxrNqRzrl9z9hH9FaT0HgaQJnwlVV
sPWoeAD9IAxdQ9kqr3bapEhlVg2tFPxxRN/vkBatCmyLH0TKSLLh6AxaypRVyNJaTNNVXz6X7ZGF
5QKiLewJseTbI4HL1PSSdh9yMzfdQENR6WSblZkAQlm8wSPh/L45dxWLcX/nbyZU0b7C+owRya2Y
+J0Uk1irjnMy/WrichohF+NozJ58c4bFoBnbGKL+LH3QGlD6MHzHyq62+3Cq9aB7wD3/JSHObOpd
0CVN9Fklhm7Fm1PnfbqH7gBZcAIYyof0yssbAK6oI4LpxoRx0ZCYzBm9A59n1HvW8vtQ+jPxxpi6
fReIkihYHdbTnqNl8LAKERcM3HddoIlGi63Mgqb4wJLz94MwTqFnh7Zm+eiUSkiPY61Pu+7U2xTX
YM04fTny9FSez68myR7YlBWjfM/aLlboqmGC20hcuw312UisZEzZeplejQZ5DqMReQH90f/le1X5
+F4tyKw65liqHsgkdhHoMhIb3CwuUmkrLu5uMfJJ2l+C7uLSpnlgn7YSYCK1Spn3JxYZ13DRxSoi
ek4crXYjmH+VNdaobJnPEo6zlY6hfweyhmL8GmCu5q6AcLvXUqCXuvkuVzMu3qDzfCngybUauArc
kCRwRNG7roeslcLNrZM8qoRS0PZ6WVuJSZDZHA18HcbZDd8zskwyj4UcPJ+SQpCBwd+Uymrw6vww
8PjxA1YOXFJ/5nEyh34t6yMnvVic7lJjZiY+ZZlyzo2EKm6b5J1Tie53eIXbHD87aTlpzNH5vprA
FVCizHySb9kR2KDyWJoC7yIjD8yN42eGtxbAKYq0J0cvSSBtyGngRZh1MJexu/1SaYDZZdgfck6F
l7gPNiolzEE3JECpzYd9wpnMhgWalGCphiI0GjQccfgIg8aLgC0mZy7uqK29wID3xwLaKip/TUEl
1QcsYHnqggpazf0NYkOeQp0b+wQ+j6n7JspGt2VcCrYCG2VR5TWl2B537IDxRp7guCTHZHddA+zU
XLvhydIGwYeSVmDUoEQNMZUXhY65nUYUAlUF/YWXl8TXJVYczVr6wYZ1Cy27TTVOBBGiOnpiMuSB
tfq46Nc9816mO5O+LRUncSqf5igr9b1v+0VGEgNhUVxNxxvyZAfNmoqmYQBulRbeQiQfdcKds4Ss
/JMJGexUUf9dagVnq6h9mn+A46t3k8QHI3UkBJAeq524XOHmcCkOhJ7F5977DyoKzNKTKU+ZhXPt
OFKfNLuD7zYarxvKVbm3DuN0CPS4DResJ0spGYQ0r36nic0Q6vvLqu0eyOeipcASjYZwBMAz2uoA
yqGXVmCMxjKXZ+2te3At+16qTyr/9QurzttGgi+zMN6cTrL8trAdJFCoUvaC5ZnLdtj4IM5xIpfo
6zzREVSa4lUPdj1HusD0KdZPp3AkkK+pRmRzB4zKUhs5YetRaSWJJFfI+0p+tOeAS6B3oXj6/cgI
6L4pZalnVAMsaLra/ZusRRUHe647pKLZNLAIR7ok75jmJhgRdUSsv9Hd0pdvwbMpRxKvGMWtCDMZ
hoaWI6ZYIk1DwOpxe3Gbnbntcr14NRJBaY6kTbyEFneewIA0PZO4Eb+psqb3xZAawjnP6OrY8Kuj
GPGr8EKmV70i2T7hsbkE9J5EDqUwfwt9zwSHur9Z3ZC9fKkzxcilyWttN9x1gjDjYAAbQJQHRe9/
cf7iyI3FRb6x0pciDubMuUDHktapPnuKq7q412k0PtRlN8IITUyvBi9xR7nkMcPnkkWY0m1aQl22
zHFGvPiZ003tTgdU6nDgW1CAwk/79NwZkrqMQCxwzPKV1WyNrpoeDuX+OJkhrLKO5cCv+e+1MAwB
AiICwMa5sawBoZUvULSCpShANotnYYGBp1qZB02u1YNrma2ClaPvow49hy2bBzGoLQu96GKLuWIx
xobNIUWLhQPPNcKF59E/Ztw9d7xvVJ/JibkMWZiRKoeSJyeoC8TRWbeTOgeGQL7J15JNPNbd2XJx
fm7FgBJj17P0VUwmnrJR78V5rxEk8O90g4cBn0ZNqBsaE3pLRTeUuTIcZlASMvb7jUfrrMdNVHpL
sb0bVVgx1MrBfKwt3xN70zox3gcnGMutgid/KK+3OpQEEa+YOjyzRjV7IZGjcVfSSfDg5g/3oMIJ
iuKPHm/gZbE3ukUoQ8GM1OzaluWlKdSerNo5P4XYGAX2CdJVa1uPoZuvNuMrjaXWHyfjWe3FfNsA
YJyjEiT1Vkwr2LyYf26lrttPbDWRUux3rFTG6uuYfJmINNWuZFau2D2mQP5o2Mu6V4zy0+lsJ+Ve
sM6dhe/m85TDIRpeYK646cvl5i3VdiS8UL8SVhwNudpb0Vcx6lJ/rKsee9rYm+pIczfW1UnFZ9ly
+ilDtuXbIQL+4gZxfVdgTPGfDWRuX120r07DMbTRpZri6HQqE1ATrrXG+ibXCq5yxNKHppuXLVA/
DZZmvaGf9Jg/NU3ecSZMnX1++saeWFd60EPlGdCK8Rh1Wq0Pic7Zc9KZbLLr1WXDThHKl/yPxFZ0
BGeowPmzVKoKS0cx7cUllQot1aOO1m9cIMt+f7gnfObYs3ptVJQs1IMDMJWSl9G2pHWOL/5zjusF
MvgkPKIOVD1Zyf8rRXIh8tPDnuTSeny14daRZMPpkKWZDXSaa4BZGEZjcDSUa0YQtM5iow6HWVRB
nU35C/CteBe4XY6dJ89BS7WKtlBB6VUGCEwcrC7/JaLB4B/iEEW/nRCB8l2VL9Qk+C68KiivK+vn
YNs9V7ymTJhi1KzUUHWp7UmHPyXh4sa4dUvyF51N57vNC0TEqvqd3qHwQ9CqWko1JsxmDP5fOmpx
wD5c+HCR6v00g0+G5hi5kMGDyWAClLQeY7zmEFc7g24V8YS9CsDxT3obnmF0teKSzY3SRCu1bvpz
ounlOuXyVfspLcBczSc3J76eFSBT+Wukd8our7RGFNQEznoYD4wQyybaFdUwkkZt/obGKie0HKkH
/w50VXlRqlZ3UaUCOETy2tYnlMvUeFCt7wqtKpwIWLHA2CRl3IddLIBleheFtAP6X8rHIjwJvmEO
r+fQi2hNSKd5NTotqZ++yRBDeoPx2qAUsrqT01c6oJYgyfwNcHagAFdVKain3wwxOvVTlhjRGDwu
kZsyMMj2+Kry5QWtna/+O/8Qo0sZ8hwV0NeJ3u96SCYSf7nMIqpCrbKWoRDqof1y7OOU6Hwskwus
d0Wf2U6mjOGKU5mUE/AZT9gQgBfcoSJBvBYIrmsz1bien7GVjFBI8UtVcgWZlI+cba1IBIO2Za3K
Ec7nS0B11fgpnYKuhEotEwcUl2yH1WdtaE9u3j3bO2xGZVEPcrGNgQZ2LxI41YVS35mz7g1kvh7O
/tS/yrEGHrriaosEpPJ3fnWpU/5WvCNt9x38djk60iwJGqxI+yIBH/pje7dDV3klSm6jDOQyaoXE
YZhqvUB2tmR6hZINf/7L9nfg8WPKNmkYg5wILW4aP9LmH9wuPBWHL7meWrCP2BZ9uF+wCdW12hC1
Ump+kiy4KevLTmoO3yQ86a1IGJ8yJ49iSRZiuiyQeOSTqmfyEiO2bo+k8IQze1vc9TbzFRQ+qzOm
knzaAVh5CcFNGB9YUYnXc85vYv3OWUVBkzsOE+kmMMkSMY9IOHPLqQnqqWwC+Qg2GxiXzKk7abxN
8wIlRYM0nU70NYVbQNCp7ypHMt8Iw9F8/5pHK10/ccIbXYjk/QA+Lk6mYRW3bxp3OiQmRokN9CbJ
xzKd/q/IVuOLMQZLiGrqAKL6Sl3uzoBHiZ+BNHu93A96RQZzNp3olykFZ1jfrQeOZv4NhYpc6AYm
0qG5tyEXO7nHeL+xUUfzs2hRMjRcadbYKbeGf5an6KDifo8lA6Bs2nA3NAhurVBLApKNOEpOugNf
NL0LtX8SeaCaOPf+rBqkA07j0SuKqUs6u6QBHjtiRFiqvt6ta+teR0VvP1lgRpxeoSfwSON6699Y
5hTa/gDW71d0UM8DXQVroGAr+9ASqYT7lSZgrqz6MyyRxQ4cAbH0unsp8f53z07xSihgAq9PHyL9
zkOJ4qbZlqH636h3ny6x1b8llkVjW4bwsdVRTzWQSTYpfU7kPBFmHJ+rrc3TwFiErdQD2Uu3cdnh
Ze1iqPsOqw3nXhYiGtrKAi41fBSqm439eo5NErbknEZjG+TloLaO2t1Ukpv39h31PIc0Ol5EnXNG
sIEB6MvSQtRv+cmnUcq8bwXB93T11uxgM7sxSqdlPh3ZrVO+MPmj3HDy7s0wab3mi0jYBKg5Fgak
sUxjuCTfA1sQ+Fffr1kFFZ3LOu4l8zW5vfEtNqKLkec00NRR/rf/nRAHIKXaBg0grfV+rklvE9zX
Gh2/eekAVv7pqVYfz3n79/+ikK1JIKv+Cvs2gROHpcWucDfpJg6LJfnGwKcMQSxIPs9ThTII7tYJ
2TLuZRpRXFUwSq0f+iNJu2iE0BoKwREqoIdI/zGjIWzp66gdbwiZfSvSMmOrG7Q0pU5IcHxDSZtt
oOERdslCfL1knWO0TQO0497Mm0Tg1Dr0aZq9nK2wYkTYE2lCtC33qospFV740J9BI6ub/Ixxixur
YiqmK25ZxI0uOPF7mjcg2hv03NFf4MhnE4aJnqXgYpfT6wrBOEdaPJfUwBMCoCeOzcnkOqpIoi4J
8tuYLNYCx6BRFUguFbHLf91CKP1FzZb7LsJjE9NV1VUPfZSex7+OmFaDsfpXRawVtCQhXmuLfFT7
/FlAirJefdsOuW/xj+kxUrlsQJBg2kCtRnAFQ5Hec344Ei07Aj19bwG1hmt9580elGAjuLJoEI93
XiO2KSUL0Hl4nJDcwCM/44ctacMRD+tiAcZF4xLZ9xR3JIs8gCioSGDpC98SJIOncg7zSlTEO1Td
BOKx1KKBwpJmJLtz8pvsd1IMBRvo1yv75G6tC11/A7ljysSdO0nv4QIRFUMDFWrFEnjs8KbhVilK
Nnu8+inMhzUHU62KFinLIFF53EuJiujXbStiBYO9+5A8nXoBcnVG/p/obyMbOiGwkpEJH3ZAcsGt
2NnxNPxLMWthGrPEWJ8lU4qIhoB6OOYv1/bpiOqT5ZiTjUo14bd9lb5adIvRHSc1SlwMxcTSPRMu
POwa6Fb6g86T3icYwFhW9kq6s6UVU5L6YU4CTWSqnLFf9g1xlondqLnF6uk5CLbK+hwmYxxDt8ea
hNISqh4sb08ttK/sdZSRF1rD9TC8RXBC+bGLmNM1CQpL30Eu9S8Bpc/UuNly4pg1DUJ0CWo2cBob
UKnsksDmCS2hFh/yQ20ptggAAyQbtY8/n+j/aWxPXaN02ucKaSbN331e26ILwcepYuxotSMVg3nv
NHketJ4FZkQ5omc8k98UYCSdIfrGnwnbU5cqIhqtCMhO+zBOTqG6lcqlagU3X05IoI3R5W+KqyvO
wgpBw95Op7FIvgzycxboxckLzpOGUm14xP0n97SAep2ESTRQe5+ZrltyjdsT8t9uDMy6uSstCMOW
Ggp384ATBMXf4O75SZix/Nk/tYgyBTPKSPnLRTmT6Og7pTqCD+yheNr62VGcYSjKOmWrJ795Kiiz
IGumzfTQQG2shOjHFTmD5OKPaW6OGzQWj6iSyF9T3e5IKUDJYkX6mr2eoulmPeO7nYWM73nQYWDd
I8Q90TZHcXRBL772rea1UJycjFsqqd6RfUSq+8eyqS1tU1AncRSJ/fucRbhIEiwKisDHqdezSiH5
9hUVTtMwYZzNaTEon7jMqB+XqPQaq9Wko5ge3wJdAFhVykYCI7jayCBC33ZJUqOMwrX8VSPun4Ha
HR+fmnFThvSPSxgwUVsPiefYXJgTBJBFDPnahXFNjxpB8ayvUtCW+6N/wZrPqB1vU5Ag25eiC5Ug
EymlFPVsBTWsrRCh+CqFfJUR7n+aZf9y5noYZKqpxm2QMSNEcq01rG8Sk5LGmOOTeB722PBy5Clp
KGGWhF8UrnjyW+niLe1Djzu8GOrWPlDxNeOEgjtMpRSbrXgEhbHJ5gn2XvJVTPnECybk2qcw297o
xT1ciKIoNfOUBmKMcf3sBiqzRLOaNftbCSDs5FKOEQevL0xAobDJuXkPZSwiOa+ZhJJsDuzBxLeI
SQXGM5ojrkNrj5MFIFYizH/SLaPTLuMVeIEYRXBty8K/59qJ70GhXHkyDhOPSGhuAGaIJ5FBjr+W
GixR50G+wgFqtUz2ZTevQ1nmCg/a+WqfRUmMoQd+GvVxIMnydoDKt67ne3bn//wi46g6ug4MObAq
vz++BzE9t4A+q7rwga7M7WNAIo1YXVH572PLjAfPxX/zW5xhX91boTK7Zojtsm6YuFD4cZar7U2/
poHng1CWsdH+kJKRvIdo7k0DsbobCx2myJ4ugfRNRRCuP4FRmA4LwOLcbaJLXebtvUaQhwshwvHD
S6jBsmQ3JxYRX/ZTmzMF6rvSmWulmb+hKqUi4tREuoZBCJwG1xuSTGNLBetaCeUpBM5q7jWJder1
rSr/epz9nuK30isDDqMrflc6V3FQ1J5VFi9zNBVXNweCQLjjuh3EruQynFynKEoYUZJF0OMOjNZD
icMYzU2Pwm3/lngKYTiVu2Ad+LUpikb4deHrF3LEN21ErlrZPPqKY1u8nqRsv8DsvilmQfc0On4F
MFO8ugl98wCZxPKF5tovn90ph7JuiJH+ApKScXWQ+803GqKvT12D7h7y9Vs+uCGx7hdbhYXQaTdX
t+Z4FAuso51Wm+bAK7O6Df2Ua3r26VXUw5MM4eGKj/Tf9aiNH3ib8iWsKC7pnARTlGBLaRyplf6L
6qXH3D1dgmuwlHmNqc1FjsPAmREFJj+gPtaUgru52Uy3EeYkoGUBdBU6wcgdrNvuVkW6CdIjM22n
YAktvRfXkA05okunj05Vj4rVBkfAsteiPedYPlaOD3rRWZ2ea3PKJ/exghAirrPCFolP1nyk1Qm3
8Y6WDH7zc+myVqRdrGdsdeN6IeQ8c7iDPJ5dcO2+ON+QbU0fZK1v58D+q3LwH4G59VnUDSIhw86V
tQeNaZbmExzJ4ke4VkqI77+YQrrsjuJnTcr5xCQdRwiPk/6wReK15Uq7DToOn8E+9QnvO8x83wt+
jsrlYu8g+0uumhGpc8he/gp6JGSexBdhUJ4EP6qQSVJZeKyHvqeag2PIPHCQKpuPwaDuZQbR8Lf0
WzP00dsCEzTDZMi5t5QKhwOOYWcrpeD2VNGubmdC4WDeg+6CB+Oozz1uEGWLWQ5FV4vJ0T9zieKU
4T4JS9N8s/nMtj1d55VyCW6DiYY+cBlkmKkHDXjQYo8iIrxaSzFIvwJbELoSdiPrB1eTL9D9uPYp
wUN2UTFeMIfO/YQjAQP/70txmY81WMSUb9aW1VfrxNVSyGcBAmoAtRRBp9L2cC7ojFuVu0fczV+c
9OmUCMRscZ7y4l6Ex8fl6q0N30aqZQbndCZHld2zrJaEbGY3Z8Q/us8KRwjuQkqxyqw0qiU1bzNV
1MdOr+uY7XevPJ4Ae/458ZBeC45eprTtf1nhOKMSsFvjvCjyWzoyXDNAaUU64IEjcoFRFW9XifI+
KZngu8Af2cU3VBE36hewgGVkK7Wz1UmXTUwH+QQLuLk7HjkfK9DArq7FXy2FVX8hTyglyPl60c/F
3gPOwVwU61XsdL4Hm4nUVDsM0eRCB3WhslXY5tF/1Ua306P3UGT43UhLmlHhDHDwgYQbXhbEfI/m
jz6Lz9j3HtvnR++m8iwksCFr9CBBlDAqco1LTp//P6AtsOVxW6A5Gif1CFR58Ru3aiai9YtpV+VM
WnZUi2lu59OhYXk5tYDlQo/PZFTtPO0ppbSZ/wgxr4+WSenVWYZSBGFLGqKRreUC98pDJ42axl1H
Ftp3hFw9G/dnXFC7JwpdjaU3ZXryIQOiZxDn54TSUHv9STz1CxIjmMMcgMPtpVKsPGL5AMX2n4Cy
ncVIwYbadsIXP0A6I9epm+prkbAOcG80S4kn6rOOIaFPd6eAGErBIsLp6HM5MnzA83x9p8Yhv3wi
MvaYuEjpHxRuEp3fOwFhmcQ1PUgGThz3Fy9XftMKzYhZHkHLWdoxPggVuuytBwwgG9d9PF56thft
+/bE0wdiO3DRsNDiRs9uIueoepvItHroKkLhqwbRS28qKyGTJr/5kPmzp8rZEFNFeDqjHUalIeph
tiughQ0oDH+8fDYKqL1Gn6P/E/EqKgS+yr3mgcKpVvXam9cJ59lB+tIb5q7afXVQw9VWr2bLTycI
IS/hgtqXR7Ac+zfSQFaIJggtAnJle+dHOepf09EtI2lV01MXQHAzY0D0SHkhO+/Sk7lgtVgNd3cB
Dpqe2nyPlUiSY85mvGHanopjOtpq8rjzgVgFkybCNEZBV41GkuuIwD3BV6T9xTj96Kw/Vy8kN1Ky
h0aXCvQbKkzHCe3b7O8Bi8pIcN+jns+RA3WlHABeM8NEx1IlDRwSTBbm9AhRHKQ3BvbchscMhHxz
338FAQPmzp/+hxmdZ361e9/IZSKFYaxMKXIoQtMRTIyIxdj5okoqQJTF3b6ZpzagbzsUnt/8KyWq
p4tgKG314R1NPc27GJ7nEUvn/NxCndWzOltTp6l8g3QDmWZPksYPj5UTYAGxpjHuLGWDkylSvo9Y
qmJAO5akTgJAfKUYfU/EvN9J4D2sYUIdI8ue7ZIchVzJjV2xNkGuO3mdY5WknjAPdqtomz6s63xx
BUEvwWLFuWHqYjaJ7HvWjJzuCnrCkMwg2dsN6kBIYr1NCKHlvGLkOxyUP64aKVCnqegB3YrW7QyP
tRhSMZOyaIcGMCN2Fijtvfpr5RkdZL5TwfsA51CpXL3JqOmb1B+BcqNA4kQ1WcSyszhuWukw7E/K
7bmHrkw827OOIRQUsI/w9mvbMyjWILGwoZ8djJJxL8d0e6ga/A1Irp5w3B7Hdr/KxaQ5LhNSnhWq
oNGEgFVq3xgWl/NhCFK7o6xEABjctkFvO5+Q6rfLzQ10f3lFzIb7erIreT2ejxjF8yGylChUQu8r
sXDIcVg9M+r6B8PMqNk+m+NwrF22lKBmZOihBOAE1ttKeup8EK9HNjxhPlxvpuBhavzqsoQLCwLy
xXK/7y5aSQNMXfBs+rmumekLKJ8+P6ABTvhqjWZrTip0WpMlJ/YSXdcjhvk4MiIhuyXSnixNH0db
bD0ncoOwlRH9ARggJcIrTQS28tCEIGGSCSg1SrLusJ0Yoi3N/TCZeUOhshZfWIW6sAtFWYhI+c4u
zeUbWKs93KbzCkOubw62UP6SeBTLFTM/Xy+7hftRXIVODmNkIpt5R9+gVvjz7EreJn1CStH1I2oA
FytMDBAYSVaYK1pQ5rvaLH1w+IpGDjAal+lxW1Fxtgi4NzXtUHKzo8B+6gWbNrO9669HErvyMwxX
wo2CpyVLknP7s6hbBGH9egO0iV7mNTv2K8JJhskMQ11LPsR3D9TAT2Bnxi3x4ZullhU2L2DdxwSX
7SbPHoGjvJUvdt5HMNYG4G6wm9NjSYuLKJHQu+5dAwrXx57bQC+lOHlkhu7YaW38E1+iYPj6IJHr
mhEhyaouaJnJdDBEtfRm7hazL6VD6an66lmmOs7Edfov1ewwe2kAoTqMYC7J+QeRwIeUBILoYUBC
9jdGwUjOxAZ/eaKTcFxwrhDCp8UB7qqu3FntI31tB8Hd2SnbV6BRyBOYNyHfz6l2tWtMrBfxE9Ut
zEwoeAQP9XjBUx+ecetSuAb2VgVZGiWhpHs8k5g8o7YOu/fwnaoUQjgKjhXkSAq6q+4IytYKQFF+
BS3d93eNsGvZ1ogQg9yQ9trylEbwBuUgTc2vEmUuHRAukStBVkQUvTb2S9PUGIrMOwCvBQ7b+rlg
EnEpU4lrKyNDeV4j8xmBEh0ppprNQA5qWeYkVsmXAebVO+HVcC3DM/p0sgLczcvqYngzeskZ2pKw
Vw+2Oecg1grfugSU+Sp9i5ZGiBRL60vtOZ7sa7FSBt94u8Nhrz6GS21JOF+jF5/h8dTwxS8RqUXc
7Nl5CtlQEgSK5kE4lmC0VNaEDkT+WSArjRto6DnREzej0wijSeYbuCBik5a3A9UVV86DmLII+Z+Z
HBjvOeCEikGMclRpqtBr4zIW+/QKAEAxNyC6GOAYme54CSYqxNtESNomeBhExjYZPV206vD+agkm
xKmt6SEodx/IQAmpMstSLnKg3UiQuB0559kpE0f/3y7KI3gX4zzm4tpvzqfVVhOycDHar06llCTS
qNWhWj0a3bNpSEVhbfAusrenSWbvaZ1TAqDMriIsjY3XuBeOn4G4OCEd+yw/InuqP3tVCBQtsoXM
XQFtfwDUhdYIkqw3Eay7E4SdgkD7QuQeh2R3nyab+7WNCIlV8zx80HkFtxA39ZXJOfDXnc0piPjh
pT/BkmaykIb/bX6Ea1nXd1JuFeqIwK8cgRTNjamaIxeoAs7ZQSXlAQo53t7lpnFmd4PzNrdbnGHx
m9Kb6CSexqAGERiE/bgBQydjCcG225FwN0aFA3qVqMzcVnD+UX7Dx6hS7xpjphVYryhd+vUcAn5z
XEoRDDTH2nVm9HDPgCPXLRwemLqM5nm5/1ninE64mCZkL9Xsa1C7QZ5PBVWSfTatjWkNcYcj/4a0
2LVdWLu+K/FxT4EUOcLkGowo592dVqFqFvXNIu/S/6kEqz3Hwjrz6l9kROEGkj3E+DnHrmat5QHz
tWxU6Pnjzd7pq5ghU3IJ9vmiQooqi8KcN/JmEXHx51WbfcUydUmcF9caJCGeq24QyhWqYoYGUzCz
LsV3WRqmNKBSQi4n0rMtLc4o18DeGim5qgvlNI3A4gssFpEkPN96747hXYj6eOo7owtlnZ7K0ohd
6e7TiYSW/Ki9CPSQyD27X2nrnMEZFuOBSa+ssysDqp5omj2Mk3gXLpqd60PgzV2rEtLYRc+lirSA
ylcj6/kaagpFmpll3OmXaM2A+1kY4bFiXFavGFd1eSdqf391BIdQBS5trx/byuqDjyLrJiYsHr/r
5brmJnV3L6t5OhB/od4pLeoQTyXCIcnyoQWN0zXLxunqdXAgOSaPL2mlbpxjNWIFeBxGOv0Nn+YI
dFiWO0YEcVFaD+nwRPUE4TIZxxxPrVjynD9I2T/IXfHj/2TJfM+BPwyXPdjjpEka89V6J/ai/z76
VviZTBlqnNXpncxPjPb7NIjYXbMlQp980An006LztsIbw22xkrh2n3f1aQDsO8wNM7ZLDDcS/YGG
21Jq9EUNHYZueh93/C+XyQyue8xDuxiD8urYBkDPsF13C5NavZADMfPFsSylyq+ETEBhx+AX8GbS
jXWH3KAm02EPikApbdRKq+NboUPZGr9QSzURUyVmCg0vw1S62A0/M1p8c5vDfCt15VnFrBQxUkts
akMcRenCocs780u65EY9lyMj6MOt4X6i7cRycEWv4/pFANtgdJN3hKEGf5jkVoemLrfffZmW+L6h
TTppnpO0dgldvvIEUUhqoA/vJH0Ouqr6hH0hGeaePZsBf9Z0EUWQdHbRk3maPgvSxENE84S3Bwg+
ydsy5RFqNRmPLE3IJKxW+Z/OAJuYRyU9zhX3vG3e9DkHrP5tOa2tO4DLapzKhBVmCoDDQgNxeMGm
WYSUsv4Yxo8pUL0ZkdoXQ+tIZYah+xq2dJvuJmXWBpFGqo+PHPVj6K/6bR+znffz9hjXGW7wSrsb
R0vREzEGxjolQFlkNomlssKXX6yn2MTJLPTyXSQWjS6aYuhAZSlDWx79gZvWH7T1qAH4hbgLq56M
obwfVVRvmjUh7CzA5LeO8Z5xDJWviRa1nXzeOQ1Y8vD3fzLhot/VKGi3FFg7BZRvzd8upKfWLrB/
qgAEoeyTHnLMHJDXDfQh2Iz7tL4vmz38nmTbfhMhaCWScy767tAiw2krUuS8Z3HEzBCkMSUH8alg
eW/R8R1q3TcRqkULP5TEWN7bOD/T4xVPRz5eIUxy92KvASScHt1suzPTtgd1IaZvUfmmyQDlp1kD
eWVMbiDYGBIylo7RdvkBStj6QhHr37753CeEJqXx4TphayU8kD0xN3tUxo97zh+G3sJclcdY/2SY
aIHOu+MIWJfnxePVqwMhxM+rDICRqdH8Iu10i5ixtyHstBZM1x6+THM9Q6umWcnLtxaFJW3KDDC6
prZkL5xhbsQ7FI2uP1vozr/KE6Da3B9F5kR2zeqdqi9vtbD6CKKnGgLkZX4PQRMO3/JdL8AH0pCq
o3o/9IEWPOSI8S6L+J/H2s0ZfoigeGTwaYmfFIYKjpRVsZf63sBgG8l2b8JsNldr3GsZLdXfPLOU
UG/kYeJys2lZMDjQRIjkJFF/8mBP5XJcT2SsqN98k7ll9zzbC0NnjCr7xrHsFrfRay3PAQQG/GOq
eCVAlH47H/3U0tY5TGBXVouTontIkiJv2n2JaWKgKzoMpMN94k24dT9X/8r7qg6ItB7WJh/chIXx
ZHpVxh9dnXImSSAiiG1PEdpt7gCctMs7bp68AnxKQbCO7YMOJ30Z5oZoK6QyLz+781yyiwqrzdYZ
IdjoEIIsM+ORTN7OLHcDZf0WKrFPFv3Ecm1FvSFdyG/UFXH9+JRBIo6GEFEpd/z6DRbqPNeg+Y3F
v2Yg5vX9bu8AYcvuFeetz7Iz0VXh8lY+7UZvpo9fZQLUPtF7hQbyahE6hrJxFL0UTbgeK0z82rFS
UyPf8z32ETvGK5wgyh+FoLuvui3OWjJie1/F3nNJwzcM3YPjn9y+mnuibbKO+FjURUDVg7rhk5/n
emKQ4+9OA9JcpvSf4MX3kE4lfwtJfnhtTnxp/VmDtAQ8i6a1+LjvYx49WU/M+6b7Dvc5ymr+zFm2
EYFW+zjWtGHS8GzLt9x/9kHZ1mCzfy/Ph0Tk0b4h7LtnJHaMcLglxbNQigOZ6S1lKTZlur/3Wn9A
+QmzOqzn63qaaBxnK77L40nshPqbCb47jdYFLMqH9NYIpf3K8ENg7SPEsCit3HvadaEJNu1tsDAF
TmPCn6yQ+1Hao5K97l70Z6pEYgA3xpMaPTruFhwm5GDIAegQXz0XXLPxvowPfKSVfF2G7fb+zDG7
Pd7DPIjdnGevz3hMV9TW5n7wZag7OR3vR5q3vBn4GS5VOWyRqdFMObn95YNQljlkG6GreRobGuLo
AR/JglqSlIxu7EGmBfmsqPfGYFmO+mtEATvKNiVoLz/vibhR7D1IbF3hZaYUWXBvjnfbVFgUL2b6
iiZKXVI9cYYmBlyI3cNCX7ozQTKgTOvyxJN8/LycP64YAwUpz7pNWwTq072Cy06XDBc69f03iYyu
EUxB4aKVbijep455GqCuu7xaxPUbmC15YhJaDJY+LiIT4FP4TdX1VGRm+6KAkHk/+Rlee9RHRw29
xI5dkvanW/MbW3/ca52riuwXnMtXbVFT33q1/LvxCAdgMNgO/JHfZgOm31GQ4YR80b2cN6uxgLTj
Il2U92n6M4dde8xzvhWcXQYhpGa2gEYsntxNrmpkDd5gr/k0amXxYWnBssK4RFaqK8gpuxKUK44X
7giZCRSuOhkN8A+nJyLITHVM9Tqx1YnzrjDj9ChrqZl2CJjQOREsJXW5WK7Di745BInK4sCq6XZ+
MMREKl1oq1CbaLJFbUUvHRBmT1nOu4kEWq8Q+9xAeojU/JbLE3N9v0oBzVxqZ2sTt4aksjD1g55f
3CgF3xFtQ7oWoDbOEzBk/+1uGodH2RmLloELSgFLpZSbWKJil/WBo8PuJQ6JXf/Qmz2DF4t+8wd7
92oULaovWAOFm1wQ0iCIm97XzsS4lUhi0qDyk/ao51vscqoJI3fCN/sjTQ9WQ6WRiVby8r1Qbk7s
o+uYbDbrr9zBIi0jJyiz0XlNWho6oZaqoXcTOk/FtxDOQFYkg+H3ITUtLrB0foC5NrAmx2+DFg0p
sEhf3AIIDReDNHE3uertBB3zsFZkqOKfxkCkrE9YzP58kKPiPAx2OsDRN/KqcR92imrvTTmie/lb
26AigwmItv7a5d5Y2zppW4sfpEgwb1wZ3lc/KqPjVj/BfLogBdpvgLi4vcqESGUMNed6Q3BDBaE1
e18oa6OcMQKvS3+MGlrhBtcunyT3o0H8z8nDFsxnOMUZUjKh58f9hEmg9gCdoXZaopbm3YHsmUKC
APwlElWP+7pf2WsUGTmx3sij7//vkLXasW8A0UkP2ZmNmGrC/V09kNahLGRiDuPy6Th0qk9WjItg
V7mslmtU0WtQVfFX0taS1Q09bbMXyUcV0XQlR+C4JkRyBOOonAfXEraXNhNS+sWD4AaqLGPsUz0q
Qfc870se0xu6+R9OUxMV78Kc04/ZcaGgtBtOUdfP1x7uVDEH6OCXI+/Pjx/hNhNbhyZ84DsyDVEB
L4ivgoM0crDsZzTkHJLVhwlmVXMOcH/UuW9frgBRYU0M0z15lM+eSMIG2+b5MI+8CR4R0Cvz1NKn
fqjaPkNtuSe5Oq3ihg6G1e0NeakF4BPhvg4IyJoD59AtQ/ucJbTlszN1Fh8YiiKkD2rhI9SyzOg2
7pyfiC7IyBMyrIyOVp8Ov5njt6QzTf5e02Mu/KAPhSz/wMbExcY36DfuzzZXolKjptjRGz6b8tsG
y3yjmc3D2sfjGx93LRHmKKMK5qUrG/Nhbr3L2SoWwR/Ngqy/1NwwDp6YpMlb/ustzxWNsARk3Owd
LdMcrZPCgdOwV9N3e00HE8hvMn95zV29FH2u8T5LyYQllDCnc64+v5PvMXReIIOAIrv1HTBgY0qb
n/lkUcYd1OceiZZfPfEUzk6VZutBeOxGCSTBPzbCBMlOQLqHIjUjl7gNQpI+FV+ZCFfYJNetIawN
Zc8+Hpt+8CaVJpbAsHcn8SZsROFiyNy3mV4bzawCZa+11TWpqBlNP4rVfblSRUvKZ4H4OwoeNUWJ
/2IglAm+dOgtl7Fsiy20ClhlCiynbIUE+miRoDF4cCWcXsPMHJHdbdR18439+y10qSokBeZ9jPC1
qQvVmRi4TvzbfD4HXZq981vFIIpX6ky0H5ib6Iq/8eVOONpNggPZgsSXBJRt9gS49BLVE2CH3FB6
leaJZYt2jBXtJquQTIDOUz4VlAujtb5qVT6aYyoSSBlSkt6tKJQAWHP1vM7VQAKHU6JrsSGQ2uiR
UU88ZS+bzhy+fO/ym+JUDx6rIwaxTo77lM2q2zFPTG/PNaUBXliFBa0FmOEK+X/cr+TUs/GEfUpJ
M9sUnCizUg4Hrbrf7fBvEypETH4nANPZXOoQFHbnedz6nxfiQvfyjWryRJEwHYnWHCzYCVsn5agc
WsPwYLrk6/0rvrWdTmiskxE7ekhBgI8SHnidYKLX1tamiZyduRQwN+YywHol9/eRx1jJ1Op2V2HX
E/CQQNQUyhfhx7d03KGzZEaDDyhhwBtc0P9uwQcY+dzr7oJkGzj9ES2BpZMMNU5Uf5MXWPZfAxY/
8AIapDnBX37tZJvG3TB/4baXhdZWWfGGLVtG1czAZHVPlMhh4yG1p2T5MfJhuVmbKMFv0xp71k4x
/Y7iuX5Mj7cmghRMT0bMju5aRJcOO4mW9I66J9Q5PkDN8+JsKxAWvmTNdj017cB7J+ZIn/ozI5dC
NCkWhYu7rRei8wui1OZvMiOrHO0VCFKX6sa9oW/V68NjR25bzURAcMYaHi9lRLx+j5nw/9crXKOC
kM2xgBN6hp0uFeB80eNKSLolOZokONW/hSwsZ2BRUuN/dc+9KTo1VQRyrm8Q+7wjsThoK/tmPhV4
wecrrx2s6B787ulnS7tkgCe2+shUwjUcICMcm7WCr7twPQctIktEO0q9ZRxcBYrqtGeqGjGc+kSr
CxVWrewlPrCGEmVjcGmSn4NBChM4Xc7vgxZ2A3rFVxmshPpQRdnLaYc3P/x4zic47rBkbl5AKG+Z
5VqK4sVC3BSB4n6UaYREN6WncFB5A5m+YXyFHrb4/9ho1GUGVg0hkR2vOt2b0xdk3pAC2WQRugoj
rDLnNbUdGzx773IRd16hZdyqwdrZhCICgav/4oG0H+vhURSA3J/gQz8B0bupn+2iV1V2ar4H/lyk
uD3mvy2MpeZPpUf8azJaYaEETO6yTvgWRddFDRWC9xMNROOk1E6ZteMpD8iXkZc+Tf9F/3E5uuse
Ed54F08b+MMjHpUoTIe2felN7vu1g4VGnCHPRcIjTTZc0PXCU2EUSCUNJ49K1oEEMuJK8BDN5H+Q
uDBbWxkfS+PtelaLZxChT0qcMXLPYWssxMnmyiFMUakxg8pHJXBx40UtN1eNRPTu3xZEGXyf17fg
h9ACpGQlRg/2/veDuzBfayx8xcWmm6kRqxysyqsVclGMKADPHYOjnEP2+qDSONd92M2JQwCp10Zz
Q1ukQCeXsdF0qnDaKblYS6OjFUds6ouwyIG7tK4pkxRMSzGK4zBGXUM7pvcsWWp9ggdUw8vwD9K1
6kIXykKhugulfLxAELIqE8sCs/c/JCLIR2EeFTj/H5jHe2o4Kj+WQXgFGlJE7pE9Gk13GL9y2VOH
Te/zkPdVtl8mPyyZm7gmwXbr/iGjGCxjfVQXxRwrBtumgFCnCZczAmi/1LTyRoM5lsVoNefUXKob
QtYiXwFM3yrBNe8NyzwZAqg1obHByaEP7SrkmVpSAGmsPpS0pRhw9XasxvyCQ7oyI7LjhNmABqx5
9ZtUePnWY5w4SQ4mGTCwBypBYvNcH1M4IvLGE8qlY+p/yQotajE7lMSS+nyQkunAf9f0Tz1AmVfg
XHbVZ9ekMdKn3aQqVxlzyLDMABDEJEEI9xetey8vgWfuL6NEUKM1TZvr41fL1lnkoZ3yBbp4/Mpm
Wxk22DfmgXVaxpERWzJrP1xsZ4SkDPy3+AaeDFtW2pjhhsk79R94R/+oKmmzRzhFEnv5JcbB1WuI
pfFzoY9SBCqr1cB8geNqe36luKaVSSCStHSHNbO7PcfANOOUXsNtt6N2Ex5+PNUwDOxj49a94xLr
w7AAIXILWQVTisYsMeVZ2mFjjncOl8BkQ0Cn8/DFWrivBUX3p2xNVmoejQHXlUwUNjTQN79JV2g7
gH3n7Jx7EehJ8mwtZ+vx9z1L49VpLVEGBhh6wwVciUPIKQtW2xDGQ+tRVT4kA9RDEjiaupXFRRxA
bLAh3HW9N1I/hUqRjLvBdgkTzYs3VxvpWvK6r2iC07MG4iokR8VGSFKuGp4jqLet5pzCjyZUFKaj
KjpitG6L8pufw8HPdlxNP2J6ZNdWTaM+qpLGlRpn/4dapFXqjzEaaqIpcWdMkAi4wEeJDPon8gHI
aD38NRzhJtVtMuxvzMsYGUOdoJZtJeW/yO8hTpbVeCBjcF/V4+RCslg8VMJprFXENLYW8KGogNvm
/dRgkCivrOnzQBl4HDtQ73XWRx7dQwNSrwEuZ4O0x0DGzflKjmgfVjpMj75AjSYlZuYCYgjJ7PzN
hkmsItIo9/eGFxcmFtASPRySqMjrwyKqMd0q90tI8JvsO9m1AUL0sswrwcRwd/2XIO4L3wcjPVHp
r2IPK+pGIHHmp8raehHQi+4NL0pyjkk68xWRi9Fs86n9uO3cWTFXaMlJdOEHIlwEx7uJQvCimocd
5/vCjsb1CLHIi9rDlW/a/dTS7+32vQxgAXi7FlHL0xkQh6/rz9Gqq/pzM96E0LULx/jn2t/vq54/
KXXCPUy7qNC4CXRoFDQffukpcww27W0SfUMdbN5QzRuo9A7ZVPs2hqInkstdCt1xKL05qW7nrWyz
rkxizQgrsKDLGeNE2V2jR8sFhPNb014A/aHPEJxDBelMIhi937S/CPTmXQxIZ+GVSM8eU4axkeGD
T5EEW/drjDMI1mijAshPoeujFqwA6r8sqQqxvtDs1UsOQFzv3xmtqSzhl35FakRBS8JV6YQoqpmT
xqhbo1FTQYnLIV77fZ6TQHARp5MTclzwgEnI7DIwZOWDm5MeNG8ziQRvrfexrBvFVVKRTorPociO
4i9CyOhXcjWsJu8uV6OZYNqZVnby8Ykq5xhkq/gHba5sdn4dHIaR+j6kQTDNRX4yo8Z55GfYyfBM
+5KHpEugguQpN6iNjWCcU8mLpuoHVbpVbRAnJvhmOTXcH1d/6DJH5YsGE8dnxqcmlvCepJR0YG6R
83IJjt0C+5Q1dThdO2OgOrtcsEDqyptwZMMFqcu70x82aZG33yK/8y57o37rb6Z9A/Z0YKEodIp2
7bmMtF0/fdNPE35c+dnoguCYlOzh/3UXa/kRvrru8F5x+s/DycnbhH3H237pnK6cEZah9lgTtAKm
ZTX2Ch11YDEVRQcrq0Q8FE5r4BBf7zuHLeMSaUVQQC6gpNHrwaK8lzcnb/OocEF5kCkywgySw8LY
ZXV5RRTZV5AHVwe9l3OnCDFeJMIFciy/mRD1WpcV6cWwqIoAHX3JS0gkPMTShrfZjtOGGVW55XXt
PkEBa7TLN6+hWcnQIAOllDNgFb+ldXnmKDMITkPUljg+y019RZ31jzmxF+yVuPPVgQz65Kk8pBDg
ZYj2F1+Tv0Ox+2HH2UsScv0l2z8A6yVbrrQMajj0E2LE9l/Tjw2m+tolLFLM1YSdk7EUcgli0Toy
8IxJJTOXTm0ebZ1wNmJLjkQk3P4/y8QKP1KmN4lRtoXAofYhwcdHGEHUMjUfww5aWwMERk3rwtfK
PcTIirY+DZuvmpHpsk3dTFkAXy6N3wkI/DB8my7wgSAR/VZxzium6/N0kqfB4Z2Oa02koMBGOrHs
k9gAt2YD187Outi0hd27/plVg+w2hoxq8Wh4wHRUCYSKxJUjyowRI6POO7ty4sGwtg0p13gHgzYQ
B8j2GF6l9j3KbdfY9faMgwfXsAuqQTVOEVlspNxUxGddbi3u9Z9L8Ic/ag0kwmsozDD+dpGBVAtN
BySAInEuxyMoj7NFkkckxAXLRDMe4u/5lmSqXPjVpIve1hf1sjBG6lUP/ILHzRyTSY//F6qX1i2h
H8HLjDBFYzP+Wb9chhhiX15gPhSONZUv4ZrBrOqML2hNUjimtJZcHAvxWTQyieqRTeKzSfCmaOiq
FHPERnY2+ctb/6ORi4wzrMiO1bdNNBbqCFezSbSobwO/IS+vSiu2yHcN6WgSX+zsVzY+O9/DbHo/
UAfA6aUUN6PfHg8+f9e3sIlV3n39zqtCVVwzd1PJt+Zo23m+6Z7jCUZLczOBDtxnFjMOe21mH/RK
UPYLoZDIKhaZ0dRyyXyzFjmm8JgFut3tJckoju/BI02vcTBNmRC/qq9b12oMuoHjnZR0A+jevpMD
4I5WoK6dXkvXtGgI42B+/vpzqdHz5NYWQJfE9zCZ7H2RhpzeMGA/zLoOfRKwQbIkmFSGMVLMSm6q
hyAI4KEW2o8ZxvH3yYCqSuX2v5wYYHVlTnS4RZuEmgBtqVfSJdZjqFhA0LriKZsjDAtHQQEnMlAN
0+Uzf53A5pjQzX5wxDySTiW8e0S/Q/iJsC2kfKqxkbqDdBwt28ZVXKUO7icuOi53pNhTUfAn4C/k
Im7f52ODmYyEnAiMGUQe7+J4bdsgr9eRPIrAJphx6doBxkhdQx3ZxmuLLb/3fafVlaZbG6FNvr29
jMw+C6WXM4l92JdFEowbKhmCjlpDo0n+v78jAguD68SY3hzRAZua9zq9jQgL7UoauylN4MF2vzQu
IK/tjRBOILdDGTVpu4Mo+8c3j4jHDA8nk+cgYZBbLPWXi3E9KwPHmgZZWen2UGX1/Ljt2K6rqUjj
RYhwYbdGGqzDTpCdSdZCaikfptyVBjEomYAAC+t7G3mIoa+A1F1QB7taHpyz90FHdOnUe5tqqC4K
TOMuuE5wVymGXiHgiytB4wFlwQhZna9r8/cAtA/AGzncSxEGvLi7vajvZHfSWBxh5lpT8V7bsXi0
A34aabvX0FFHE0rKB3xkaAGdYG9G4Wd1LPGODYYQSKDhuggc085SEXv2W6w9Ralu0ZqgJkMQ4VJB
tqC3f1xv+QjYzrS4p5RoG8vm82AuwSGVluxg6zz7naSujL8k+sdB9Hy3poyHAbBuTjtZSEa8FsGu
1qkyGZjUFGxwGL9amZSvloZiGbPbLlM9Bx7H5V/C0RaG3r3cjpNRalJyvFVXQA2oRO+8lajdmLv9
tY+GIqKcOd/iWNxFQqOYzX3OOCR5ecs8VgVI0d+TDeQZf3x/AgpTPh5Qty66DyYsN3ZDmoeKhuUE
544nlUvX5VM7PeJsOaJI+lnQHwOXNAIUSapNRbMLtaB0/mYK3A70xAsWhbBi62/2lPoxi64CW6+o
9xUZzpVUTfxB910Oeg1MjGFq4gw9bKoHRhHCH1XA4Ub9h+mJ9ltODenQSjD94Cv09WNRxmcE9oM2
pwXOawXqzsrriAC1Sf0EaUzonrCJSM3ns+oYEuSkSuurZdZ3e3+Wd73LUULYzOv6NldLwO2t30XU
2pV3NRIC2/cvtHDOHq7GOLwkfDwO4dsNZsvRGOgj5xckqNGQhCuabLFe1uRVa3IrrZWqXhNpX5Ca
47DsP4DfYfSCH53Cdr2y6AadQIgoIS4nryEmpzn1RQLkNrCASVrAiu7YKTs1CU9+tzIhW7pYaxJg
DCGyC2gDaFALd+jrFU1mBYsbxSwRXHZueltnnCiUlQhYb5TTyE5SQA5bHAVhY9ht4g4gXIa9xqnA
Mdk1p5Zvea6ZR+AEywei82Sjc9AgSlW2NIQHAZsAqj2/I7xlTCFldJD4xHEfLmkhgslATBVrxnop
XAGBQbMJRMbFTUW682DJ2itgzfr7SkXF3DnuRG3WcrY+3/7BZaW3OYnqWCLP3T2FCsYDj9uABww/
pRu71GYQwEL5cgRrJOAz4Nu9bPfNGAbK6d37EpEH1jmwztCjXPVWPziUb28P3ZlpQK/L7tpeZGv5
XX9u3/9/FuYU466wE22uDwHvliiHBgn0TEtoFGdusvnSCfh4zLuhuYRzQnzntj2G1Abh/4gFCurv
uHtgSEfS0SINmPRNOzucpdI1+Hx3WW1Hq58biYgYrbuzMKq1iuf677jHHL94+QgONbHxAinvzWVe
uvPOUSHlKAFGmF4SFSohsxtBMcaixkkna2cMaEKE8YOqcoMQV2nC5CKMIp1DpdU8ICrPR919MjOh
7gTGOBGqmwdIEeAYBdd3aU0GwtQssoTGQFtzlMK4B+thycz4IQoHjgPYwUoD9NVq/+YKLr/uqzVp
cBioRAtHf4s5RmZCo/BxiQfXPnPlgkjgvVkXtaIzHlZsEqxO7w1mfZF+9Kz+xbnH0YQ/uAUzcZSE
Tr4RlRbiCUMzOxtrisibiOMI36CwJ3XVx7xAOrg3gpFs2qfEIvk+bBUWVIoMRUtEIZE1dxaiYnyH
pw2L0B1tLlwytIdMmfdk59xsPt8E4Ypyz+/iyYSX5v3tCyBB+tb0T6jLHaXcJBBV8Z1tysqPL3Ze
TH8wTw4VYTSElXWzt/FRgVytxoPejtbm3ZPdMgJSOvx9jaG/yLBSdNi4oDDQadel/uav8kGwK5Y5
Ydi6oYqge/uygJ6ZJuMcE3w6c5Az8sckWFlLoNiZQBy/QILWLfBGv+yutc7O3KwfI3NTfnufVNyY
FSNGmgp0/55HZwXf7JhoJggR8cVTgEdsMxmD8NEBDyKrstUrlEoxnCxgEiga9NJwNvKYqUJnB7IJ
6wzQsMwSnsXomTuV3QYlrbjOODjTAXzLf1jsR3TmJ6gRaNoLlOCsYuwME7s0FF3T6/ik1g106I9q
c6eF0MO/AAyWRUWrwFUY5yoz0wjuj16LUGOarP5JFpohyxWXApQLGQiC6Fs4Jd6vfJoQxhZNTFwc
cnEQ0Ij2qZI9AnGFmc8AegsbZ8yPOeYnXWwWKPx2EuF/6bkkU7FjgSmyLTO9KhYU8obksAMhCMJR
uvDTE59KLvJ1JUhCoCQdUBJccXFgkxwZ7dbJOAc+KdCLZnBdQF1aNMaCb/pWVPMVzHHGV/omqbEH
oBVfpzWwmvbxsfwKkM4zgVnaHO3PSX4K1UuyerURntpcSyfwmkDcT5NQ1vZvIVsZq2c4nTz68Hqa
MzcfmGYEXiU0Pnn1s5VQKUTwuy69OUjOAx4Zf+AkqPm+yCrXz7g2btfsHWokUIpf/ZuCS37Y+Hs+
IwcfboixR92v97fFOodM1YkcEkqB6lMEJAZglLgZtYJdhOX4sQ3Kj7T4oziIDQvZtM/GHHT+4q0v
jyIQSfFXJH6IA0WAiWZyHcC9rLE6Z3/Pfwc+cSVqX+ld6KnuHMsn++8fgg0Ka3o103UMDiQ6jRuR
ysCyQahDD5c2akqsSr+xr/tgRBl+rX5oCBSrKu1SJ/QK4y+dCcwBPbevdqhyzrEHcp8nzw+iuk+o
vh1lBpAluZgKRyFufG9Xofh7Pz2JBXg/c8ys5zKIwSND76OE+iXjawSkxdiNp5K1NadbiNRNR7VH
XSkTslnppL9Uw5IPutJD0t3NWDyX34U22FCpYtVn/bteIWyAPIMXVrFZ1d0nQx0BZmotWal8XJE6
S/0aIki+ES6ZJDh9VuwTy1SBGfewHAiSxRkJrV5tF2N2s27xb+nvAR4YqEQtBqzVslJlEAklbYuE
CnrTuuQVhnHS9t8IRh44Je3bBqofLk+ESwl6/Iz4BAGtnbO3G3ZX5l/GXRWyuKF8cszrC1/85/Fa
beDq9sXXxWWbdTP38Yrgp22TcQLB43LZlIXbAu3T84tn60gWhC2Ji850SVv8W5ChumMPJzpxK0BN
UE2HgDn7bRhgarfPRxVvQASSgTibuKB9TagzpfnN0eIbnl1LhhbwShrA+embFBkkF6SjwaIDJTg1
8icTIQcHyaU1Ha1P89Yd5SI3UDazVVmxj2HhM3jkMngMhto8J+fMj/q6j5kx73rlrBs/GdMGA1Ev
pof3xRy8l5uZygayGskCk8Ak7UPE+8bBXJgvxjcgJ4FyRu+cA74Uhh7qwWel3mOZOGfyNmBwV3Oi
UYb2q2FeX+k46KgUPbP1b7rpBA8A0WcoI4ZdtrkrZej/0L+NkZB/cJUko98ohlExViuDcxYWBTng
hpfbl5UmY/9MoW+9O/R7GVKndwRmAuEwitBJX8eWEz+bxlf1bkYupIgBNTa+1e63ymSylUW/aBpk
Yi6O0x6fHpjgvkTa+l0Dv6M1jDR85gQcS4Q8LBj4XTb2oazVARlBBeb7YVgxXiNg4YWnIUgjt6Go
6MSeEKdUeSFUp1S9pFwD8aEvprBORoMwal82RicniiFnHZuGbU6o8UIZJxkORR2RbYay3+zp7R+x
hL9zENthfC+g0zNA6gr73JhriogSFz7JkrcwlohJ4g8kow6hloOizrLqVRvHZrN6Q5YIIuwP2Teh
ElHyBelmMMimxMDhwABC0q6JdntNgdN52vPnzMr466DxWzpytJbBzwtc3xGcTmo41iq1AR04xywK
otY3tRuq5fokYUKEvUTARYGCoR3VFmoYRbnv7vG/iCRHHmoMi0/zoWZQlalkfoPEYs2eJ+rZdXnX
prlvWjCR197q2fNEHyRJRwwrfmH2m10f6+etQYrsJuZQ+se4DDAZDs1/w+d4qp0U846q6Lx2hFNc
l3Os+5cDZOOZwmZWf+L0FELURVeKdLA+Lk2DvWOPttRKN3FIpj8Dt+SfagDxIe4NZQ3sBRosW74o
asWCS2sPdom/NEU5E7mhdYSG/0A5fSlHnXrHHVNj9k7tPfkiXLbrm43RGhkfct4BVqgknyUb7qLz
No9FrqEW/GKZXPMuW3KQ9qcbvwPoKKfiM59NLBLmn3ytba8u9HuNRSXOc9TM8LjJLCekpoXHfm7x
goBB1cEDcBIXyussuVKhEyHXH2tBHZbp1pVJaeB3+1uDRr99p/Lh3yeRCcd5NNUOcF/CrMDQRXXq
8R5TxzvhReZpg9pOy+81sZz+qIIR39PEfnFRFcx1Sixw/Twh1JqP8czhTheYFK9QuMrhJorfNssA
V9q0d4mciUCnK5yX0bpnR0WbOu0I9+oF8TFTyK/zunKSKyKbtuvpT4yHB2negUGtw4RoPhn/Prv7
a4ObDoyA/lPtYggSwiYvER0wj6HPEidhLgu2xHkCsDduUHgh+lkXXZWkb8QIPJyo6tIThjkm0Yuc
DG9faFLjRaRVmvB26Bx66bDjB5SDKVxmUlguehLd0RHdN48p7Lkv8Ra6HxUEMpGIfL08HnOOeNtP
qA0/abXx2AzZnWLpDoas+lhWDdPXdi8+LVN5ZhoJOiit6dIw+G8OYoCwBUoqWvNyk4gE86VwM6tg
RllUyeMDyxZKei29/Ii8FuN+XPhvEbKWFjyhXbxwkOfHNwDH+suSD8erOEHyDwdAeswfDhovfocv
emstlaczrxWIWKmrGIn6zto3AhSUaH0j5U6yHGcW5vJpnv8B/GSeYmjlQe3lOl8wTcqDIOh2YtVQ
vyQPKNIM8J7QjPkn1hu1O8+DcDWvxZl+xlI75XoCwYX0aHPB0N8gJMGi4MPt5KjORGSpWiz7qdT9
UUsG2AagKqkrML4yeCS2pBfE4VRTLfmGms4k+4ViQcjCja78Sca3TzxWHVySfnP2QQZtVfi1JjfP
h30ivjq71qcoy4NdPpKsoYPG3Lg5C2WIZnnRhxrf7Np3zZ6TZbpgOlbC3aqTzcX19JHlwiy2PyTB
11ltcJyUog8NkRLvbHCk6mN18vve/TIQ41YHtq5VBMztxV3MsED63tUjVqvYx3nGqgEGml2/s3c1
TpbTvjYF5gzVapFUa7hjtwoknenDNNkqmlOXVyMpq/BGUB6zsA2G/G/sX7/V7kagZxO1vcJlBQDy
HTqzU4S9REf/FC/XSrwpMtH2Fqe6frD7/cAq2y9fyOr0xAh3YgaG8Nq+HH1h/zJj11+1Y7lvJUo8
LZVCnuGcuB2yf+rgu3+bDGiqG6Bs9dbM9TCvIMKVWNf/u7PErp+vaQ4tZy3iX+AftRgsq9/HW0Iy
WzWqOnCr1nB9aoYJMXoEFUrJHz+khYMMKHFr3h7iNaHys/3tNK0grhPoYAUx4Va7ukLu16deuJ7m
M+5cAVMCUMEDeqff0iaYPOVB3SjuH6qK8vHRyXj0IYfO19YX+r6td4xUgUQRU6MK2YCNYskD/zJy
M/H7zDrJeBaxK2FWBDpOuVuRNvZCLdAv0Zm+V6GlaUGyrt5ihzjOFmL8XDThQN2HtVZyu6haE2KL
R0kQeCz5MxQHACyzLZh29XY7FmGmkHJfNLV875/iQB0nAnayXuSWbxrPwaeeL5SusKmQwsku4hDF
scQ6FfqT8JN4Ht04/hedUrIVaGMf5q27hcKqQEfnh45lJJP/46oL5a3fiMwhy8zwrDFerZbJ9ghk
gXxveh6qj/Qo9Pk3ivjBViCy+hqP7U3T3bwU0o72zGwA7mJVA5IqwS13uIY7qretrdqZ2K5fZe02
59OUvSYW5PJsHmbv8gewp9DJItJ85eAV61XJbVmF5QUqslZoOq2g3k3M4pdiwINpDHRvoJWjzuib
RUY64m0KWi7XCZAIDPI1atYap4HejFbStj5G70Up40654w5Tm75B+v1OsSBOpcr2F4G7pf2K8amw
cUuw2OnpojiZExCCm/olNd7KGYELMWXvj/r4TrgmDqebWkmgaP7rH38EfCQnUd31Qdksfm9bHq15
Y5UASjVsC3nrijOxtGO8veM6vUNWNJRaStT2009Lu2G86XMgMDKL5ZUo2gaWU32VfnxkLyfoMmcT
l5tqMZuytUE5yj273vs83XejLdfm4owZ/vOyv8FiKdErFcSiHSnaFJv98MDvt03odEsLp08/DtxR
s2oxGqIzMUepjk0y6VPi9qgBX58wFS6+sxs6dwHLf6VZx0GnJ5BTVsBr98wDhneqwku61aozwQrb
fAmAhhKlBaV/wwnRJKIS4h21c6jHrk99mZ0UL5ABoTrAUsS1vKTV4hCgbvNnNOzYlp7W1T0aWygG
NphDwFdeFIUJp2MZgipxLn+NmAJOIOkOlXGAv3sqeVw2b4kjx5TosI1S7k3y6VUULEMW6DJ1y5EV
zVEcKcFDSVnrkciRQIm5GOj+GFyWMmOPEHehN+l1XTDKk8Tbi8xgp5osUdKUCLicz+x54nOCHlL/
kh/D9HswTarw1yVPKXHAi1RAoniXzjVm/6hY2LLaR7fGcegTSfU2RSyvxr47iC71kExPQmK7mGCL
RSf8fnIEfp1wOSXBtTFRxTvuh00CXWsY3cE6Zdof4nbLxmsVHdjGWgTikvHH6ucy37HdNKQEm1K/
ptiFUtaI6pzna5eRLxPmO9zk3Ki3ntcBReab+ZAqvv/x3PgEk5obyAnivCFGDiLRjA213yU5CUPv
KT5+FPk5smz5G90aQhsn6kzmtA3SZaezQK+3VI6xgSqEoSNZNKIQZuHkFKui/e9tgMfrA2m7UXGF
L1uCLIOgYMi1vYVlwjKGrz6ZX77W52QyajjXJ3G2Lw5mA6lJJJTaUg2ueUkjBg5NV2iTcNjbA79p
brBoPaAYT7+a3L8UoqaCpL/JlIPZ3IOXcx+YNl0ZRx1hTLEZVKlM/NMsrFOJSleNk3oued3gHrTy
/7XQ2PTaLTmN0sYBFaHgbYXadj9o2om9bVJmFVBzMgKOS7BG9vkS5QghsVrtQh05sbA4VN2RIZS5
UuudtdL7cPTfneoL4zGe4dbSX9sp8iGo4UOV4ef2uylqCpu5weVo6MI0Z9H6HZljvFmxZaiNT5yZ
U+WjktJkfmOVPgG88O9afriSdJ/NjS8gzP/XzEB3Ro5dsI8zS8RCCYMUV1Fo9MJCnfugrr5AfsCh
rxhSc+se5oFvLGHOa9VwC5MzUWba6uTs+RqLWEMhu72Xbk3zlgTsydzcJdTDtJnfzrqCG503OvYg
5lKyqhivFkRzOPXPG0952ppxImTBBlLZjlM/3FARC46X362ZlcvsFLrtvd6XaC1wWvILBrb69HGO
WIQd3CsfoS3aAgzX9CRwvOceR8zpS8uVTrmBq6GJVNSXvmLvi2Q4+Um9oWifb27tNDCMfrm4QJ8k
NBdy0nJPR8MrTfsqNkcTNB88sunn5DvqE9CFKFXKqUwVFzjlp8NF/5ObnYGEhUUFJpJZD14pdpVM
aY32/5HUEvCmvejDhnr5EvogFVYPNTuBMVEScDBM5XbFIZBWPYWry2wBuFLWNhy0pw1LRwI7fvKq
PoVoQlHjLGZyiJ7ercg5nVRMXeJg6/ubwGP+7vvRwt6LC7zhrP0txVCPOn7F14MuM5+NVoLxDDJT
cO8JqSv48/OVHliSL5fl2FsVcaL1rY+68oDM9LOaJWLQW2bb8wG/2bb3pVbNVojxnjFG8238wYO2
ryg9heBoDwIyXXdMSONZvfkfxAYDrznqjurfYC00bpQvC5Zg6P03JfDH5bc5CjQaMcmBxFk8dYjZ
uXR69fFx87Mx9+mSdB30ew2naMy0FggRKwYAFZ5qg5D5NY7uSOXVLSkS9sIp0IZBVF9ffMYkmDr7
D7WW9zd1zWbpw6He0H4yK6Nv/vExiONv7qxr1oSBahp+RS/y83ht+oYzxxjs1zN8BBe4i5+660YX
0gfJXqsOxxxNikJTRvsCaEhWKMjIcCXYDKfgp7AFCvq5XPFPHYyi3fn2TUO86qSDqBCSFWcl0d7h
KnvRBgB/bB24U7YEPf83IiddZEhUPUQKekoVNL3SMjQz1cTWx/go+FSQ0glE6fD0RFH1DyXVGIlh
zWm20f0N1H29XS9kImRdxm7vo1rIIkY7k7AOBTYiQXGgq9h7hWdtGHaRMoAXIwbP7vN93uCr5ArR
lwAtkCCcVG+0iLvC5MuanaPMMGNv7cuwoGgoTu5c8Tfv0c76jej5f02vq/9ewkPwKZfTTukeO3mr
Wa0aqDsq0ttMw14Khk+wy3dPFNSNiqA/RV3Olfgzr7WUnqm5jkK3YEGBWgIwoA72EUoNW3APWMND
90AuKh9fLLW+tIpgkD9drcCK5btDq8gMxjNOus0TaV41wvTzGks40ZQew0Nm6mULk8M+Qx8bXrbK
eDx1nTEtyj6MU8CA0SIbXdHg22gXLytk5gGiZtGd88711SzMp2Z6gKwlkznS4WKJnwR8LkpCm/HS
WjYgV96zgtS647R6luuzHSJk0l9be0iNfc4mb7nR9/fIViQed9HgdzrjsGFUzIGqDy6A1vmc6Bth
SKQet6L0drji4jP6VJ/rWFO4m1aW1zlRIHF8L8B2TMt5fYZ351Poo/ofRQ+qd5HEyeIACmD7fkTm
zRkn4o9/dgiK4NGnSa25V7pCLu2BFzp9uIdxZp1rjcZOKCQAVisiAwDeHbkKQ1ASlyvOSfHvnpty
4Ke8Ife1OCqAVCUpy/2Y4HcH5NXWg6leIoO9xHj+KZBE80Tobw4iEXFPsE31pvCD5GCy2P3WvxLO
66Srhd2yUmKMBbyEhIIANhqLgRQ7FRf9y9seukq+51MQdR4IbNWMFbthI02Okd/GHlH1BgQlxAxP
gyHYProDvuC/D85+9WuZFkwQPe30nAyeJV7OFHwMMserYA9sJVraOSLoiXMj0o77xTC8wAJDce8J
4S+LzMc+9q81lfd1DwX90slp0a3s6kyHksr464ORJUmxaKDSut+vXAyVGhdNXIsRMT5u+AVN6gkY
gNrm3b8w2wVWOqrG3MAVYeV4a84+QzuEa3vs2mcZvAJRZPuLKgatayqziIPOffGVtVfzZyoLu+1p
dDHa1CDuoS3a8CwSQXCv2i+UcfFddDCw1hVucJMeiJ16LBVUlsA3y+OJnQS45vEhd+cLPqiS1EN/
dBk7dGLWJPF7skXfWgUbUKNPyXYs5wqC836/eA0aKljUMokpP8u75X38+RcVdp04l0T8qNerFyJA
FNx6PIT38pvMuK+Z24zL8iST1jcKWxHQYmCyv/b/hvc8ylZbh4e4rDOnh6LhC+QIKUNdDY9pR4zq
ODvCB3P/YQTtOR26IC5NMAyap4MMXZlnBX+3n4sbFqnZjUl2zF5pnitovUe9ypVRW015qERfDQIp
33RtAz5cTLgBsw9cMpJCpmp5gZVlkz0TGU5Rrvi3GGHDG/7px6S3FeM7/8XU0KsdvnvnarUG+/V/
ghPmO/ai80++AX/7se56CpjEoAb6hUZlK+8858k6wN5aH26kO4fxwr77Dvz5XhFEBDgXhT7+ttBI
/I6u0r80pEyER85rNVecG1408qCzdj1Juq2xK0ncGssxoz9VxXmGj8kyopJ7DPz8CryRduOxZNr4
SrqFhFTrVNA/P6W6BpoN2v0txC7VYWH6NLEonUy7Sq2O+YeI5Fkpo9hnoOsR3LPB+x3KwFZtLFWI
eH9WRHwJILJvMMlnnUXzV0F4rS+6wRxJZOQ9SMCSRj2RdTfg4XYSazS5Uk4kmp4ZGij1QgXyoF4P
+rqVmqAO9kEnqU30RwnCPBkIkHPeDCfyIUQin5OlHWWCFwqPgKSKzz3WoWDU856ZJ8/kx0DMS0VK
sZqPGnZI4PShFJunyhTRmeVHcryM9frnOKm3GC1qIAZcRukGO1pvcplV6+q12Er+4fXcMzyhodgc
cZqO+kKXyRUJ8J00W1gzy4ge0lLtKZqaOq3bRZexZrFbK1E+4FetqhIJln0n59roFAoom/+JJ3Eh
d8NGkhYtcp0/eL6bE7DxE1Cylpsz0tX5bSVTyyByMMN0mrUCbmuoT9pbo8jWTW7iIdrcShPbx5Eq
hHAipUfCacSyTIEOl/2+YcSlslw0TJkIBHE6RkwDFev5dd/2HAiFgdtv2RxKzpZ+kEe4yBeDZasf
55d2QWv3ZQe5KT0aluyNJOFHBSdponi7upXxb2IGB/vL4wsuwPFXweT5MYpKuBO9KaGC4FMjvEMT
0UmY8hkliBAc/nRLKnKRUqllfMB+0tyvn2bIqO55CObzwk6E9oa6v6CmPn/dFBiaAbnbNGrsrg7Z
PBu9QF5TGm7RNGRhnYAs5p6+75Kdy3HqVnDktMWfm5Cq96mA2k9e00UldV2GbIJVRH5sYSXqqL8G
aNAB/sAd/ENN/1E8Ex/bWMXBWG/Z2D98+GX/u5u3EfU+hr26gxc606IX8gb4ORupESezifMQEadf
vxoWksrAzSrZQEP92Z++MpWXNWIKmDGRnyw47ZHi/lQdMDUq5OQkP7b5cZKNGSik/w04S5yRdqgF
2rDalWTDtoYlAzQ3jtBYuV5etfZb9ZPhVmjO7iAIXVaUdSOyPVewLj2TmoVIR737vXjG8y7wWPs9
M4XqJVGCg/fU6Fl9vqEBiqlWAZFfnJzpwPHOUjrPfdCC2scaQp+TQ2Ex4vf6LjhT1Od9jP4N6bJL
Ybja0VVz+KBPz4iKNxahWGlZ0c8oIR3V+NiicKb50qAliHDsDNpffNn2k+Rr5+IdRl64QoBh2v/R
6q/XFV2ZGYIF0fuuwd4wpOwrUJmiqNl/9PikLFM0NjDWQaYPdb2tkOSqcR1jUUYbuZvEZ3blISeg
ap91vNjUEoAeA56XNqYEyjieQJal8H36hKbDnMv0542Pv10AphWdzbGwwRnTWdnv7Kikkh4Fk/5M
ueQanh198f3GC5/UfGtE6UB/0SQA/CSQ8VLUzAnv08WkklXqDEPCu3LBQabTqwNaQlTvT6m1vvrW
KZOUl1Eg0vF8Y23cZ9HyGFLULq8xpV39WfnqX2IbZ4Y/xcDUMy4pnO/BFghq7+5fxkHpQ8Q/Xbe2
61y7E+2EEv+nkFmUCBY2uqHVsVBpYxZlkc6h5H94UfmaiTaeyw6IOnfoWjRM/7nKGYWdGQGPvk3x
PV/mZtL0/JXBF4ny1BNJNJn72/L65u/P+/zsoTkide9orzUNMg8tPoFUFcCOGluZNDYjBD136RX+
pEtWPNcTsLFoI/S5j1wu09TBG2vSdK8xxYIcaAuN5reOU5seeqzBILdodbLUxWBBK1+qiL/1L7Ea
MdG9T9PiOnNn4BGZL+L9nQBY7yE8/Ghelv7L/tUU3Svctro100UL8GfwdWnNnQybMKPG340VpT6N
0oVN+Odt7DVEvjcW/1aDHmcaBqKwxKgviEy6HQoWmeGlAiFEZzbwR+1cB0iwOoFR9ofIhJhAjMID
eCDhcVDIYd+q6zPKylJwqS/k8hCr5SRervoiJf3uEx5JLd1leVYymK7rjRy0tb4zUuojet5xTCmx
2cZ/u90QzMokV/LnrlehbHn8xyK1fG82RJWv9MEVNIL+2O0vlRY2atrStRRCXY3+WzPbA2ZYBwWB
bKotP92IxqxhczCjIS0Yw+7zeQQTcEEYsIVNkv7YgvPVUIg5MveuHUeCm/VidzMod6+rAQ1qrN2g
iCsWj5auFJ/4il4sgVAUwRPt+YqQypw5ccNYIcVNWCdYn6FBLhghqFdkkY66+H4Jh36gbRNbTZ1t
1SlqveIUwaEHRp85NTVRbo+eR84X+bXI0NQ0Pb1H33uWy5+C4YbuHQS9IDGrszXdvhyo92b18h+M
LSDXBiIcJxKuUmWPg/fKLWvITKSm6c4IpIJh93BeA73wsrV9WPP2C1r5my2C66YHo5sWhw9vwUcP
m+3SGvcjXwABHiV9WpKC33vJltnMg5GOB4QEbkHXOeED8jj2OJiLHkBa1HcUUu3a9ZNEppyzKhHe
UC45Pu32PzGH25OJRpdRb6UGrq6GFvc5kefafY6/n7cPsmErqox+52ByVFfQBES4Vx26BPWRIgHP
lCrwCybCS27v9nUyAlpdsT7fkyQ4Iqn6btD+h+PGIqaytFGnl3x2DQ/gRwrvxyLKTB8EnSneJ1NK
e9cg2xy2BOy662sfKBA0+G5iV6erbPMq09Xpjf+m4ff5ANTpFMQdSddSVVVkdyROz2Ymvvh3sOSa
EJdUQ4NbARjG83jLuJ7k6Grkuo8Ky3xft+1BV+xmq2a5S3m7m8z426KPgWVhW7CMtWvDP/s8iWbN
dTk5yTnV2wnWeZZbCugSqwC9ImLaPyh08jkm0BXyU+osjAb+TvVCv4Q8Y+29cJfPri0DSyNFh3ys
RvVqfN5vBwnuyCfn/PK8Z+yTZy6pD8RwdmLspb+DCCgGqvaWd/IXJaKjrm390wu/f47uezz0zR0U
lvUJWeA9Vzsm+hPfLAh4yOUUr39hThjVfP/OqFI+WoCK+5mcHk/grBq8AhMh5AL/qqdyf/B45ZTq
J4il/LSZCUS9+ePvZ6StSvdcNN+XlzWuxlBMsddeyaIviNeqnL9Jme4L3mLwXDpcc3yM7aa+1P0/
CCWiffaIIPTwH+zTCHb6CPQHeXFvKmGqeyZEAPEjvnSuwZXy7MkSdqGUktCMr1aD5Ii6p6Bp005b
I2p0QC6kojZCjqXRO2mouaWKSu5yvDH1JdmKFa0v0f3NAacAqgKyF+UyfX/Av0C2v6kzYVj0EgO8
yQq90AB+GX+ql4qmKqFPBjP02dTa3kA0mRUrVu98FZ+lk2ceRZ6Pay6BoLpnaE0+6cNASTSM/uXL
Fkea32KJeKXEQrfp1RsUH4MNwi31evpNmPBYCKAFJFyaBcKzgNbRK/eUHchR+o6U8Zs6sD1v+M4J
sG1mb8Qb/zVVoys8ABZhWf1U95cNpc/WvyzUKNg+8Nab/4uF2+8OedA3HB8esGLwGYaj5xGmtHcv
N/8bcdL+xtssAaFKjvY+/Pa6SDKKR6iuaz5sgehwruMFDuDidjZTH2/Cx7wQ4JPAi6LB60IUKfdv
RTN+WKkwaXcJPTkpSfJ/fbADypHj49WFSkiaevrije/DEsr+hd+1kMeTHywuycrF+c3d05AAxzC4
WT8jT/IEDNnNT2RfP2w5XTGtYIoB+H8HR3x5Q8tfD2SZeLPB3+y6ktVeFh4rSsPsaCfHEbVr7WM+
QA1w0bREmuKtQxTiZuHQ6FdM2uHYh0ndSmgm01utmhBpHUt9jUqJEPJCyzKfBxZDQctVU12JquzK
ufEVntgEWEogDMV4IzQBj+aYUP3km3FWhuFe5YYiX/DWkPM7XElhY/YWpKzsuS5PkHtOQWFrfqqi
7uMjyxWPLC+4MR7PCJrTRXqbpqWjM+y1KmJOqG9dV/phdK74HLfG7FqpV7UqsFpqsjTHj6IsMd8J
AeFQPwXJ+BP/rsa6GBz5bWH6c8adAAC712B3nzz40+3NdTdOgkDSOXdl5l6xSrmvzLP7wk5Oy6bu
n3x9EBTa6KjoI1BMxH4ChEkw9n0z7NZW5vCVEK/mmn7BQSikWM6RGQBz3CapCvme1Z+2qRFvM2w2
GQZfKTqTZnNunQvPGWcVqTCL3sv9zvzKDJeH0yJnvybpWNJAm+7FSKVbRDK8tMi2bumYYg43F0rY
BqDiNxhn5avYcuUIOvyAv3O8nm5RTfwmJvDnC5TuH+ANvMm7qnZIUJXR65XyrlKEZ5XjATblkhcA
coHrxtPTYrLYexXhoux8IelPsY6I/T2ATjHVomuHyXXnPAGWPJevQumqaBdU15Eu39/YNQJvOL2z
8V3KjSer8F9Cvs+ab/psuJ6oM85cwVyiqeUGbu28uFGWUEqPd/1/m9ndPAKEsgi3105bIS0Kp1tc
cOFbcXnm8q+OuezIbHYROp+29sEP7KlKr4WeG4G/lUpy/REL+O5mv4mBXTbySlYiUtz9jvGgQinA
vmEcQ+ZDd5YDQm20XaQOqEdQBL2GPxV22GVzPCHhWw+78zj2NscsjY9KN9ed8C0QGYEtxwKyi1zc
l/yxdZIsJd64ZsezMJy4ilg69UJb1LNIK8qj9ryceKodmiDjGkcZ5QikCa0Y40TRWoIcYQ9BAm3e
06MglVRZLxmqq+4OlY4jBd858jC6uAcEKuM+fvMsGRxRDq/FjTansE/SnGry0g4VTL2DUCs2JZKH
nTyGVKPoiYhcNfV/Umi2fYE/HznRg7y9KvbYoJCmNp1tovth3bfVfb5s7fMMDnSuQmuc1gv6aqOe
P4HQsIoHiFTpmhHM+MmHpKZpv6o7G2u2onwiV7pmltGcLJmejqSeiSTjoYPfMnPh8fiHmoNEyfwq
+CnvOxqaVtrp2mUBWREk3QXccZXG4vwiJE6a8VTmWunA2ZGxlQZtg8mPhQz4m0G0TLjyQLvwSnR+
M+tcLfNTuR7tEtQ2jDgASLbQ6hSi3XthLOq4TrQWRxgoHh8+stETWAczg/9bEIGTxrR1IVGrsQax
55iqSzYYLhwbTygk8GyxVrWvyLJT0uTxvcDJaYX41ZpStV8XoSwvB0WzLLgLZ5QkdD7dUmfr0dDM
HZuCEOob0rQnA3urXtB4YPFMhKq9wv+BOUztI0/HvPCh7p7R7HIy39Q5RPxogpuOQ5hZnSKRuVnF
3dTGzc7YKhleGe8q9gN0yvsanA9DtDbkzOF2sM5dfBjLG2BnRJuwF3y1ZYEWopXIGqk7agIAHLMW
rUHtn8WIxmLHpe2lAiEBG1EHigQjqfDBRCTYhCQOyaLyWrMnD0Y7XMEPkAYoY+6KM7lIz2GWIyNZ
6dlE8o31wMzOn+40Qyk+7skDiJzwvxwJU/Gp/uMeK4JuIbdx9Lhf0Bm5c5WGPBhdnAsCdZk0LhDm
ViSJETX5fDI4o/RAP48qsOMNEq+a6c7OSOjtP1iPEvIoHSC30/MPUjsLJT+ERUFGpPADBTmCPC8K
9Cayn571gr7M8SpuG6W9m7DM01t2xD6a4Ns/jHmmOQeHJLpZTNUE+QxSwQHTeFAN3d4TbwzIsa/w
0JlTrEinhyt9BUosazRQKiqESU0vcSxGP6Pao06OvnJAQsSGqhVAW7UmlkVHmFaUBPB4TJYrS0FY
S9AhmZv/adbAuHzfwioYOHbQG6Bk7HMd7ClGbmRzd3wQdEO5w85PFt2HoAhn+tB08iSoctLQlkgS
vhf8iQNYQXw9//DOTb0kvTTc8UeWgEASPJFfHdT2nWnlfJjFBqL7NeCCenWvmzEehHgZ5EAO+mn/
YduCxSxWnzkVJeYb6V93oMmWGBA7g2PnDAIeT7DgSAHUrA50cJbK8+H2EwFLgzrBJ7ZY7aXdlKUE
CLC869ieT/8Twhm+D43Eth1+4erL3Fxjaz3tAAMWOYAFAOhXD06jS0QY0INjNruwtoPBSElWrekS
VoXaCJY8Rrm7e6FzpkvGfwV+D7VyuH+BU3uIwsNhndyPubBo2I4CoKTrDssib+1VB8IyVSTOzXlW
mI1sbsl7Z7hs1+Tf0eqxGfQIOIOXHYmQYXK02gR9mSHr/tM7jeNTktKK6e0SUpRqPKlJltBWAyYv
Tg7ggpOJ0jQ4qh8NlUl99hwBkfHnMwY0DnKaz5xASA0wylqzOCRBOEFqAlbMxEJ/b2GIKtbdGAwm
21i8iZICNZ/MQ45TcZUehr7I6CvShKYhGMgmeAuJmeYJbzBjqwziDEV2+QfD+Zk3FsAfMRZt5KlN
nCtbpxXWojy04++w2rZ7vtHbiL8BSRZmDFE4IVCWuXh7iADikQGa8rTr+9yswuTmI6qkbeJxsD4S
OV4tGXfMWJOXSC/z8lcFMcn1UVcajrPT6OlrQP6XDWTd+FRh9JnoOp64PMhGc2Pk5MkchGJCE4Fe
GbbVVspPXypCkf9gBQVVLn07TkcAEzEsEhRKZbbbPBDmREAk2BZYg5YZ/SpI965ce4/yl1+c/som
DJBXgCBLQx1Y291U+ytzXw/e6sVq/Tepa/8dd1A8XQiBshtkNbn9bcemBfHsZciesuyVYwDVRDlw
GWJmHXNaRJ7MaR7InoB6Q/o3hx9Lzi1h2Ezkzye84s4T5NT41SO9NKB6gax2L4oFHjOoDoJmSdPw
m6GPvUerYY3Dn+waHzTF7KVlRKnKywaxB7aUmzvNXnPe41x82v6R71Va5ojqhpyrx/C8Bcc04O6x
bnxlDRCTmSZTVZ5bKb1MBiDgpTlooV1CEM7sD2FuZ0Mzu/MNJ+hghMkqYdIvYGGQ1Dr5yxDJ+/uD
LuUagd8jZ3jtfKAGKGEHPzesttVZOYqZF34DMKA6T4VYLQyT+FNTKYhU09Ce4IIHmLX3aK5fcQhi
0EuGt1FYkwvkQNgVJv4ycxeIrPm7GpjkXZAn34sOZLNAR07+Jv4KTKWv1OFhwqol4eX2d3MNcirn
RU3EBs7HyDhlPioJcce2TijjrEOsQ83sRZsxSDSaf1lr5VYpSI6r2/rMgww/R5pyoesd0yKgBEs8
mvHcrdM7Nykc611sj4EMWzt44kKYaZVcwQ4M6vFCr0Li9bYIwOO49AqdAGlgyxztdus92pleu8bS
hkILukxRqezNJ4VHeRio8QfIhfkqdSyOiR9eQopaWGDDvNuLYgZCC0sCiOC4KZOU8kr4ea+T/35O
CHIJJ4+eo5sGpaMxhBQFGn/sJqa0evTsiBq8KR7EekNeP1Ow71MADxO64yuM929Yki1L2FjuGsts
nLpOoQkQcpvFPtKeM6wZYAxtJMZyXiTq+Af1GJ552QKUw6cFhy9sNbRBiG0g6qV4MCkO8AArGJDa
eAOUmnjq0Y0fl7cxLv44UCMJvhtb5ga4bMtDagZcJd5jjNdL5vex0sjohnQtrlTSIBwyCd8wJRRd
aKAX3BPkSkMumuBjLj8lQ6Cofn5NvPOiRN9NsM2frZLPcnTX+9ZViO4ZhZ1yv0TSJ3aPnt+liAOk
GQwG8cAzbX/1U6nP790kYDcifpl/R2poEO8OLdsfT/180KiqPJIoVI929Pd5f3QLxJdqV2riKXAU
Y+AHvLWSZhw3glJKJxaNpdiF1fbhYpdCI1Uf3OgzGbcO7tUbGOXrrNJTGPa27l6JqVDXZKryu83q
2hr32/BaU4GbD2qOkj54ZHxDTiKF6x/lJZH0SIGkQarlABStYZdgeNY3Tneg5+DNgkFl4QBpeq/X
Nsoj0clWyeH4XH4bFuvSekqTxj6GBzKsRLDpu23o9vshAo3BiSu0mZbilSicreQeZShdUjrzP5WQ
ZOqr2qzdQIY2RpMA0CwwEyRbjWP7VWfE/BNo+DZ3MwyAuPrvDYDCD29UVpxaySTybzVyzwYseii4
Eg2LDyDYA2pCDabj6+KfZ6Ot+2lScBxJGxOM5W6eS/kqWamUnwjOaoy8uF8sVBCesaz5gqR2UUwB
gSr2WTejG3Vy+xK6xUyUzYAhzu6A4RP2TGAm79Qcxg1jR/iUYxkVhTs7rDTxLXqmfRg43dkcasrn
ZqA7fRN439wzeNgAXy/7ZemtmYTzuXewJBUEC/1IeW1VWUf6jjCfjEdiHvbHMU1dxRNfK1kpoMFw
Tz+//WlvSOdfnyCuBZ95rnYR65zKH/kMV+JIOLnIDhsrrihPvt1cCz4wzqyxQdU2A2fW3vCvBTXS
dxiNdWyoGy86ZbxwrAHDuftM8xeBNK4xxRgf9xTDpHBjE19TZgXRA88tYcdsjjfqzjalCqfOcgcV
M3Ds1hYJ6ZvD316TPNXRp9ZobgLqFL3eFHjPMLGFjON5PWy0lgPNArU1djixQznXhrrFdDY+/R0S
mhO+Coc0YsudwO9XedvXUgvNhLWtAEp7h3upN0XRaSZZ6hnSMif7YPwjt5nUo5h29UH8QAVGnYM2
Vl2RZW9bUd/0uqEQl3VEn8hTHf3jGmnPkIhqW4/NLF6WodyyhoxT6cMbkHearX5MYqOxpwj17gD3
xXk7oPT7SJ58OCZNPqArfORG2mRUBEWcKzfIkkqyC/a5F8sfd/WlbuRXRLrVkQMlT8GDgm9G9gw/
LI0EDPRMzzjK57Vh2ee8ztIQ0D2Fr5jlQANeutOzAn4V/dfGIiVFkrYML49WVyvrgI0Ufm+aDVAb
1CpjPfnQCwc+OEejQOw7B41p8pKdzp0rU9WoeXD+DwJ7q4b0K2NEwzwPPGbtmY8WyDKfJ0hdmoFw
3P13GOYIHDuLGiirhIjRraQLjafUh/yOWl61utJQc34fddgqzSR9IfOr9yOsTycWP7ZXP+iKDue8
X+vAtZI20MyPRz1Ljxs5TCnlBGravDpnicq1ElWd/vpbTrUj2MqgEFC25ppffR83a3QNY4mPmzXs
McaORx9IZfw4lMyC0DnhRvFPQJXxfUTM0+qBy61csvNt11+3cyDnI2ztsGkmo8KhCgJPB5Qyi/LE
3Cl7hsiY3IadvOigLcpkt4+PH7MPV8FWWeVRenW08ssN/tMMk0KxwN1tLY3H7nSWzRj1kwoI/gYl
D/u3t5luXYZYsyI8qdDBrDRzDts2HS+DGKatYrI5AmvbqNRLNvwOiNjz6udwaJzSqzEf0sxYNwfl
JaogIXhqcPqRRcvaAF09V+JNg101EI23ImYGrlEhS9p4QkytlSM6cUy4HVC6UvIpoXehB8yp77jM
bdfT03mV2w1xf51LTZgU93EJgFr8isvKNMMO46143iWTZN2aUftmXc8fyytY+YrGjw148AZK/bu3
KwFRX0ARodFpZ1fz5Z8EfcY1xTB685u8VcVMVkicvFQOUijvW7Btxg99C9CjAMBQxkfF8PXJRjTd
4uiAV2kif1JpF5Q6NZcUIS6e1rQyfBvpMnmYNoUDVIq9T0Kg2nX9mgEN4KIblrQcecaWoib6tCmu
e1WW4v6B1v8aw6J4tp3/px9pZpsMyjYnWb9iayZQ+rVWn6/gzq3HIbZov2LmGQ/rIyNy53WEBDW1
F3uvMbG7TZnMzTbhDDxJRyJLjxsUu7kwcR24V1NhYFTLSzDHdeQuk928++dz99gILMqlqhpzsqts
gwpOsM9RyqxK6gJT8orcHnsettczZBvjQeLB4ha3HPuT/OvPiwwrskWTtgYYLA9RsUDvO1lcBlnz
KAnNSnHf6vxYFGxXWo4tpyT2VbFeyMwGhyyC+jd9VpYF9SaROtm6v80Ry3N6U7wiXyDB7Cumbrm2
Iu38PJrOp5a8s75HR3oFa0zbJAbPxSie2Cusp1ZPI3cTt/LpEJkzJ9tZv4EENXisNj/GuMlQLbjk
SGwLixKV1yiXGpivHoRA5A8/Q4R4+5fBERkyhFGhAODU/X2r56c+aqcF56PAqOYrrH51/+0WE4+T
ciIefhXtsXj0F1Ef0YE7jjXJNP6XJv0z9wwExg2heF1RcNnZHnCivCe0COh0hja7KRuQQpK5TU59
RnikqSiSCFsb8lvQhb/EDeI2oN9wnqh8AK8qJdbd8TJDnQEseKYFmWMz8Fkz0CJlQA/HAHb6K+Y+
J8MhYe6HA8pC5fK5xXJyMJPEJvZOZeACNi2Ss5GJIk1BaEhXD2p8gH6YIjFlxhgoNt++YzM5e8JN
G0+DXwD9/b79FCNT4u3qEwImFqeXmXzyGWc8yncIUuxbkAPI/ca8k8P67gHez29aK1u9bx2mwOlC
wcSw3g6cfTwp8JpyjRWWW1VGRWH818U3mFfIBIuDaCHpWGUujxSsEH8QAqYBNqmcsJkAGABk6cIg
24Kq2yuBUASjtrB643S0LtvgKOqCYfn5FpFv3tssSKXsQL5m8X+yHbHbAuPyPGcVsJnWwEz67Y/e
2lJJM6HUfxGay/xvPY8Kcqm7xGeWCciWQNxIVAjPDCVU+Jtk6sbZz53Xc2HJ97TeeNiLNEkMe7F1
dR/609Ay2PWIuelOy9/Hbpa593x4e1GSNzfO1e5cM2TQSjIapVjWI24NiIpKGNfKau8xHvfi59qQ
j6Mw0I7lt4VRhQ/RMF34mRr8233M/ZiO7oRa6cYzvJPjY00a+4zmvveyJUUlxBykEGOdWzqGfwQZ
yei5tMxMdQS7R/zcBPcdHhvBRTb4RE6gKCNJN10WHE492mx74Us8X8bHKI21KmZ+xb58xQnAAWLc
b0YdrXMoG3csPyU7Fa6oRa53GZ+iPUp5Mx0lM3NEfHY0vNH20mHAz3RThBum7680D0YSIVPdEYCE
Vnko+nlNxouTmiuJQ8EmMVPHlQ38DVuA0raE1aNgs1o+2ifcrzMGngfmMV441PDUhrRhEN4G1Yz7
UohzVxhfr6q5uVem2+Gk9CLdU9qkv06uyBpJxvDG6y5I18hWxrrz7NQhRQWEYvzV7z9v688r98py
fwBxYOW6eF6VcjYbaf+GSDqi88WeWLNRYlWGADyta096KbHrz7Q0MKyN5yKdaiH1LkdraqUSSCcn
kcVpAAxOe8TbM8Zeu5xnCUYnEffXFsClSaXBeUQVmNVht6QF3mjJOXMDndawINxiePI5lwWZLBu+
jdn9XjuLaLu+W2v2z/Vzshg3rCuG1+XLVhMw2j8EdFB1ZTpTEfFBUfb8Cd7fdJL1r1hQC8zbaLzj
QebKUFK3o/MRCLSf7Yu7U7N1piQFXARAgr0oCZr24MA7Ptl+rFbxhE8Aj51eYnViqO5M/kiDK/Hr
AE+LSCF5YJ88onWKv1GdkZ64Rsd4EOo/Rsizx0bIYO1WVUHcCROI2a7aoovJmVtDuRcHbEHA7kyC
bj9ohEfd2Abc08t+Kx17FPz4vYQG4cKUorsM/+/Sc/JoembXjgaDEWbpJW3px8qss/KYaBdtCX+P
0yhYhTNI0sO3gmMrzigZOYOCzAAxmW3Vr409MDrQC1xNBdR3llbiDD0+XElw4OBlvyJ5xQHebjP6
Kg0irQfovFtDHo/+/j06yjTW1qg6rA+ZCIraFtQs+h1D0hUDjwo6IQiXBfw77c5+55k5f51BQ5JF
nCOyr4xwNJQenZ7vOS20XzKNCvwfWIX1fP3i+fduRyzaumtIY8jJQBgha/RJWRg8JdOJZvdGAIYl
/XNlJcoAxKDDf4P/rJQWMGpLpJqrvUd/KOErQLuHfd5CsmTEaqEBv1TbQ3cHUsSsQyIxMIqRCWgF
W4+eQkLZqv7CHHqzFAdyO5u8fMCC0y3esSfX7PF31bjmAR+R2SSeuwCfSqCsQzeE0RBt7PRt48IR
6ZArpqCQS48xwMT00LWMdkAlRkiFUsYfbHIJlfQowZAX8Zsy6XCFWGhBrkNSraurvC9+czRtf+Hu
2T6E7xyJpC4vlaJuNHISSKitnXOLVoqi/B07v89biFgjjICnFf9hl1Feg6b9XxB9il1YNlShYnFQ
ro7+MJRbs8jX+Fwo0yvtFFv5svMqaWq/O66CY5FmfeqpHWxUy8jVfEnFL0y9tdSDandyGvi6j0iV
GL/El9l6+8ehySk/TwMCqBJmZP2+aRNrw6i20Cg/NQ7S6Ce7B5wM0vQwXG29KTbp/JUgNjHFtu+p
Q4lbakVsIQa4vGYdU3XDoybvsi5vT5wuuiIi9vzXFI1GDOq4WfS7yK+wQvHF5GBlERwcVdAta2jQ
8h0F+Sa1F5UzzoJiZY/KW5GKVbzf8fGUt6gZoamgdzdlf69bx+e8sKyTV1AZmWOau5HRZeKlfLm8
3wO8eVJd9BdBYJibMV27FtILUuvdKN/eAQ5ol0BbQU1eN57rUXraWurAp2Hd2z3djp9HhGpT2bwy
FpYjjTxwplsC0t4QAQM5ilb3sxynny1/D7r8hO7IHZe8vgivCOLr4FW/K8SLXf/NUcZtm6xxLXQj
Y8x81ajbr896djecJrfDt/nbhaabKfxKPzlb++9EYEYWLHbMzaH8e9LJK3XbD7xTR1nxDPAuFocy
17h4umdBROKlQg2YhHLKz52KNgfMnf6Fhzx19BSMvLn4BR60+kSHaNWKskUWdlo2sbzcLSFrq48Q
2fscfn/EJo5iFWOtYlZqlbaZqlIFLcnNk7pFPTBCtoDtV9PcS+PItop9NiCZfzl1TrbKKyw//V+z
Qtxdw6M7dJmOdHo7suKmQwI/Pu2QgP9A1rxlSSZ6IRx6dO78h9ZnRfxcRJ/M5Li5ggAjWF9FQFkH
adw5V55l3nSRrX1ZGN4/p6mYxVdgFP76r+VX7pSdbyzJauB/athgeqZfCTJ61IdCnjjPQIPaqmIO
risGMA45psMiTlRnDNbUbiUURJR1DZpoZLykohNGHqdZR/2/bE7BSjgOKP5MDsi6hz+3rUwhPTyr
QkRydOEJshva0nYyJMLd5SYyItX+aIplZ8f8aI4/Q/7AW35GkMx0AFEC5GJJrfrJEu+cE0Szqm3U
6XgrLzxEb1bP1dLm2nXlSNGdBuTrPR4RMEpbf7g0atCKBYTwIi0yXz5JtQPy2zO7IjUSXkwfsS67
dQPUDRgfCs+z+ZRTeeIs6x4vSyZ8obQAXNPRadp3OJogJm5pRQglO0YntSQwAsbFtUyskht5CmF7
DUUliD2AXfyUZ4FPbBAEm6AELWx8dV/iHBrb0X8ETSazyzgkNEjjSFeSzgINF3vmdWWAcViyABlY
jakhrCvDCWzgqubG1fXnLc7xvtwAijTFFGFIK/7r6eNvJs9Vjzpqwb8PPt8gnjGDw1ZLgPQqp9B3
ZR5orLo3udeSIyLYN2QeXMZafvRxpi5xkv7o3cDis0jErV/PLVhnMIKqtslLHdFxlJAuATSfJ6S8
ItD1ZUB6woRKu7K0e/6zh3Q/UYyG9KEd4jT6mWHyTjJOd8aKWH8k75Fq5+ZdDSCY/V8Ht6wQT1CA
/u8KZj81A0ExhLb51BLo+DpqVeQxm7ksxLHmEkBEfqMSy1l1DgR//WXoc5ZobP8sLuuw3NQ4ryK9
dq0x5j8iAzqJWJMgY/QfnNQt/dfiGMrCwlkWrOpC7pnfK4ZHVwVGsKMp78MLO/TjlBXXw80Cpkde
V9hBzsPuj70gUKFWhD/oqpxCScLpI45bGuicem1FcI1p5K/LCK8Zohlom+R4d/Z/nNj1sklRIzA3
C3cjdHz73knlDZn0UwigatkYyM0bQu6eFU1Y4KbQKHb5/fR7RT1qhO2jI25z/Ksk+Cax/zf/QU+G
VC29bJqL+fzxx6zb6RIatvJ5ONK0dKNBA+1xXH4KzNVzp2nIw+JAR3KCZ3K05LOjlLgeSiZmDhhN
f6m1SGiFxf319RgbQ6mqeeOIx/jA/dRyM+SIn+23FpaGpQV8gb7cJV8kCRaNIWBJfKDUcp4YFixE
/3mnK+jQ+tTvDtZXHReN4Q4Qun4gUQFvE9XWS9aLYZq76PJHgWRVCxHjSLDGPtwUhLnH6X2XCyeT
3aP0hdatN1xAdf7Shk46mr6B2Q5huU2q2AnQIuYBpbpm3cWRFuFrpB+fhd/udU9RGko656lDG0Sp
qu2+t81D3TY7u1E222dR1kmiLnoD3cpM2pM8Cenm7Iz+p0b7OEzUafov9csGWDH8Fg9R9MmzPfii
zI7puZ0K9cHx4Y1yIMHUsQuAJKCWAJhLNdkfCmfLxk7qGhHQ3q1admiMYCfgLomT32tfHKxTl0Ac
Vm3VEHEGOLGQHTyVBCBEOuYHHz+sfFGhwZsGqvJA4VQE7m44YRyWA99hB/SE6q36IneZRUabZTYx
nFsg8gvOnHOdv4f0trLa0hKapMDyF6VdicX+L5cSmg8Gx4u0EWJqZrQk4s600CyTp5P2R0j+kqoj
bk3GUqwhUfq/UGWhxZKBxBbtCTHBj3xAcQIMKPZJaBqucxpaCjxsgO0PVDmqgKFT/McazJgFNzXZ
fdUd+/ut9QqRuvRrfC9omIX28O4jOv+CToVyZ2N1IxDFc37JUEf2StP9K7LWhDNzqzzdXkari0He
h0xe1nd2NDSS1JIJC/aamEZPbdBhKmAKIMDcc/lv4PmtdOmIb22gzqH1dBWTl17Ia376NI9TfDij
gg1k17wkpPYeFl8BTEk0x4uq8oWaxXJ/5KKORN3xeM37rPxeQMknAl7lq31nDdDWR0tAa7Gjxsj2
CFCLPQgcOjagT0wwjsN2XbqHCGDExoZ+NM9IgektBO3Rf5GUo7PLKppTUEYhxoZsQUJ6i3s7liam
lEaEehwnkdvcF8imXClK7lBzVDDuhVVJFgDMQywhwbBsfj65l9nf/wfrJurvYtJI1noHVbMvNaiO
MkLhwp5YDzm7wsPnlXUEO+3ZOsi3IgS7Yg8EzKH4u45KmAaMGkaN3N8jimbN89dJIcIX3GkGwUwy
Q8qpnbU8V/dnMh4lggLXUEIacFiVHyDEkzZygHHcDTTgnaGVu7rikWMlajGC8KLbZV42BtfxdE52
2DygNvh6OQae+RAUZ9INu2BpRbHVDFF8XtqT5MZoSPLcGMHWAOquMrwwdb+/PRBpYb/HVnAViQ2m
9WYtHMRe2iRn+MlD+XdCLQ/cgH0IvFazSoFm6C6ClQVLzv5m/T8AScDmihbGmz1UenvwfTDRtnpO
hCGvMJlJV9n+EItSzSOyzSgP9UkPvoNimuKaPijxrC/xdZ+jH3Vt8G0dYmsK09Mfr7FrsXK9e5zC
PYvKRaaTbzmdbIYzy+/l/u7gfUZIv848FCtSaUjj/WPG2KMZ377l0fYXKS0N3lG+ZarWBzA1meEk
djZiMIzN/4kMpiJI3eyMuj6BxnM3GMiSY5r8q0ySARI0yvOXZBA4s+mGokKJnpUz9rhfkZTcl09v
vDi0six0AoVLrOBVq0R2hcI9tQ4lsFTSKjw1wklH6cQIftAsehlktfLAY43cO34wjfVnAXZNcHcE
hLfzSP5f1ESDWzwhX5wschOKVSncVW5K3Sa5fpR+AeEMQs6b/g5sL9qEL6l0n4LO8WcUnkFvlPE5
7GdeSQAPnfNl+5Is6fiUmFp2cuHc3uME07+n4/2BPpkbA2WiwOX2Z9tL6zp+2/reRZPflwHHsF/U
Y5+Sc/YqMKKRV4O8Gha14L9gz3esn+im6usdeiIHGxvwhh2Ja3xaGAVS5oYJRwbiMZ4kuDrbCKJD
8r+O6Lgp9RHs44tIDZsJuSmHOVfMVaCbSX8EJz7AVFRpZ8IJZobh4FaGOmp0CCkz/O3ODbKhwL2H
dTiGhgJ1VMHGcSKljx6VSRtcesh/sy9orqLMjYcOpZFZV1VUMANHadJDqG+tdDZ7z8bw9kEfVjnk
yu/bh3eQsSjTpZxwPX2doz+Aa5w6sniCBoj+f1JeUmgTtskybgAtY2032MXWh4pYoOSrni1i6l7d
TY9nAu3ry3DIGKtAJmZYy2kMkhmcQARcac0vPugGiANt5ngiqzIKGKgOhBl3L4hQUU5U85jwOyGG
YGUWXkP8oYb63uFCqs8rewe4CJDaPTZVVCWhl5xn0g1HeVJlF0+bdCM/21DMxv4RH+8sseKFq0CE
RXjWeA4d7spevk4ROOqMRFYR3bsUCh4Lu/nF50aAg+4UGudDoRgdkNfnc5nPmm824fsXFMiG1IQf
Q47aSQQ91eqE7RzgTIsnbaVsKBKXn5hiigNPboEjtiC6UA14O/sRXZS7bbujrGyTp61I69tVdJY5
GwnWBxj+Tp3mwFUcUEYzmva8tMDSAkC6XfyZNgZeU4cbY04eZGHTf7tEwi1YzsknlzE8xYfhL3ks
OwPUpnDi4rHD5e76CLtjSz7Psm9UFgjgXY988SfheEKYtUM6lJ9mbMg1te4PR0QoDCBvQnGFgq+n
xxMKG48/kQzXKC3FWPNuM5BxchSvg/DC6cWCQMXrvKrCs4kKfpTUci9xAwQD96Lp6gY6arK+oJBh
90/QPZOn1OtFJfj6U77T5MBynuWCNBSIg2Y/xvLk+228LrhPpu2aJF8iMFj1ED1KYOG4vbONRuI+
G9FSXNYNo8jBmY5peMEivYehMlA8Y8o3XddZUJ8Ed5FcA1O3kiKgKtCLAlFc/VS5lnMRZyhLN+QL
Ra3vQytiMcfe+zZklcjSShBV+4hheUPMiEkr5cQnsLr1l7r2NeqLjZD3UwULmD3WqUwGDKIkSgFN
TjZrkYv2tFRQTASFtxvvHyJBHuh26ddVG/ZxOOknFKyHqofQyEGqmmtFjfZwOyetr//Q9fuPtw8s
Cc88SkghAKsx2wGX7BZFP2JoQLTbgrEBV1xj4deMxps1sSJ7bP0jcxD2Q8hnOuSL07Xa28CAgRQX
6D87j/flCQX1Jve1Uf7osq/j0RcQvtsufp08iTE9vQGcQHoECDdVIm0U8ZZ6K3nAHheHSw8Por7W
5EwTbjEn1zAd43WB+8QYluhaWNLr0IdkVVp0467qIn6x1Q7sAFlYnGzx7HE6/z/2KMBUUCkTGnGs
0I5QTZSgmjGBmztB9ookkmUa8tJMkUU7iy10RZTdfka9rDzCD7LmZmH2ilsyCU0gofFNt89g6Lmw
ynP0Z1Dzcgb+LAjNIhrySli2aMIms0D1a6lMOlYKg9VLRCkNZ9r/rDeyIUOdGjt2YtQu8/uDxrkd
7glWqFdp6+OGgS0LDGGi19mCS5wxJ3+tjkFhUl82Ee24utLs0bcjOIiFP8jQMW42ptl9WBREeTW1
7FM7TqDO4v6ba3YCasI0zHxPyKOQ3ms2bMji6rvZjhz+bgvbF7y1/lwVD+FCmkTYfGjAqt+GjY7x
MgeA8uX2/9iEb50djWl8lwbpczberFs3YJOl3ztpSJbMp3JG51pcnFRYwV2wxLtfv2CU2Tgej+Tx
dpX2zT4N0g2fNg1sH0ITzyR+8cTbtEX8AaBYFZOyZ5PNgJyYb32V+h+FV8rJT6BRjYF7YpmbE2qy
xUBpy9fspitcUuOlsfxirVUwvh5VJYC0DK5FFCfHxU/rTqmGgDf04zJKGw1fLTfUISiop0TmSu45
JZYwUeQVATGsl1ra14//WcGq0HJ5SmQmlEl+DzsAcf7SFufHIG9UjZTQ3NA+uj9KyS1oOLxX36Be
QJISeZF5vioPVAFn/WBEI/7kKIt21SNqWrEeNlBCh+qSssJA9RR9Ii39Ez1RAqVc6bmA3iEJu6Ve
/BIQ7mjKFzMTnobEkIEM5bXcOHV7fJRyMks8lUrrA2LSnWTaBZT8GrMOze2OwBsHjUEYlV/6/qnX
KOfzI7Dpr4lYz/tVEbpEFGMUeOi72pV/8R7T10AYtP+EZWEihZeoP2nP39LfAaHcyNv7vMeGj0hi
ANU/JaU7i3Z8pzh70QmPdXuW2ymODzwOSDK5sVT+KthYI3JdwAoHWfa3KKW3hye0tg6/KPIK6RMZ
kJZ6vVcf0AZBre2PCm3qdYIOwJQs0edd3ULAXAJ9Dc6nd12i7CkqlfkAIruRpVcuSr027GsLjcSG
Jdz7AXCEBCGjwZn6LrAIEbPbt6xrhtkTXjc4PaxWciUZ5Z2rHz9LNTpXBS/dW2c/x6nS5j/yd82d
BeTAPPTPbNkvXQE53D6YlR1aJOV3ShT2RA9eAT371RMVSdvGaTd4Ys+fU2bYtOxNWu0tdQKUrg1j
k/GInxbFQtJUl3DKjRvqFYNWkGWpZM6J9zrPcWKxXhHoYs1nRG6xaZfEYuoNUGcOwUx1Z8fzfd5I
XVGFpcv8sbIxqWcYIfaEWGDZmu9cLZ2aj3s6YgIn2cNn3udP4KrXbBGN7ejzAiMUxiIk4g+QVVMM
ry8kD4kKtpxbHTUYf5YwtvuFZ1AfsSbrjMgGbdg/QJCOhYHP7PQNMs2P1uq+xCKemKJ6mdep3/cs
IEaPhQFT240sI3xP6jt8jUqtCAoG+gt/znu7yPZClhNFEOK+jXr5CiSz+cNK9as0W2qlHrWM5RiC
/Q93IC/shKQ3QUWqO7qje3CcwoM6PKAJkxHAmsY0qc0SCrWO0PeslogTXHHfe6vr2bmnxyTIu1R0
AsFp5wAwkMkShN2OvaujrDJEVBxZUWECFcl68muRV0MlP43mvkYECOV9wJbu690ebgfU2kwUooIq
Km0WmnsictOwEKo27+n8l2FybbdrLtIYujRh+3BgKe5VAIdxxrTS6f7khOEnJg3pf3ZuVHwAhsNj
ftWPO+fP8ZeOaMWS9tu9W/dkqvvJ8boMwAWahI22fxeHflL4BrJwCEgGYQse1Rhh1qfnKU07Motd
+WtxWjP69C9Wkb+THh/VrKYfhp9QU65bqqQNUAhv6EbTKzy+bvhA/0HKVe32ySJwdFI2AvM4BCDm
+wGKq8Jf63EH5m2STSuyk76FzAWVx6bwjfbvRVrdLwTte8WLPI3gzGbQ96nP9VJ1Brhsnio2QrP4
84RLTqFNsijDFhY+zeGafiLbAZaml4OVgaKHWJSiENI0XHOS9vrPpt+o9mz85X5CZ1f/HDeAqR7C
b98BywpeYak+dtNdxhnx0rjiYC72ZoNRNmKikQqgn5A0Ct288hrNenBzjKa/vRKJhx0CHxzouARs
8WrHy1hLRZ2GgvsgzNlWQPrmkgWrWEOHoZjxXq+0BmSrypSY51LvOh0l8VedoDadFA54qTRBZPTE
fK1BBQeRpvcdW2n6CxjPZDugep6zly1ZZzS/j3T2EuZMks3dWAV66suvpHqwMwjnO8Zaj/JW09Nz
DCGy2jrbqtf14+Ov66L2y9swqlN+3U4ip8B1gxK3DyCoRFGJ8O9KXt6hOmvefgiLJ/UcDMKb1GX4
pXaAP76/NCiXkDzL0aNoVJ04tz0TZIgnIW+yyHXEefa6z6iZvr3TM2oyMeuocNlxXXE5wlOf6sv5
aD2sP3Qsyt9D2/nhXCMiZWd5ItTLZOOGGN1mb9jcq877XEAIX179LkNA5DEccujX8Ue6DJWsRTcz
KqlJTnmhBII/NVTrSBtvQTORWrquzO+TGtAKoJ8C8GT/VqhayAqYGnjtEGodYTpZVMvkqwqmaz3F
sb9S0kb4n6ltzOibe5D+mIOhx+jiGdffBwhTqHU7tzwly2aVjmJr5MHuXjmLMWqYu0Hix0w1vvJ6
b0g1+8sSoi+z7IlK0OgDSdujYfksrTF2WeyfV/uT9oMNJZ9iSwZ2hREujn1O1BgY+imjUnVVOYOF
j3BmspRndWOJX+XnBdeLyJvAX8P3z1jzJ/noRAs6iuXQcirn3cRVX1ICAOyqtrNZOh8Tg1fyVPeL
6TZIK++iE+7J0kl6Nm0kqn7rnRKQA/gRvduwf22Yv4iyjMIKGF5yucZ0Rz67SbtaiPlXH9JwVYHd
Nh02gnsV6VC5Wy8nheLi+VOWOZ32wc38rCzclANOS8aIwnEUJ2OMrzmoZw7O41BgyrOY2o/HXFG3
Usf5s94Jm9WH1y7f9waUMR/w3ffkNFSMQPak+//i3WiElxYMonE/Hulvv1yRoXC0KrfF7Y/Ce9Hz
2IZlu98/kDuTz1di122tuyWy1pDwrPBddebN7R2zoyAr4mdkjwSb1Ap8OqPPqCpFe8haqIew13HK
meMHc+hAARun36mAAtGUSR15GPmikzIg42/hhD15e1f44FfrruxvC9PEsl0av2yYDxiq52LkVYpN
fZyf34o/iSnhbONt+n/ESg+S+tnwjLAWezJfHSC57IIaswXbvlxfYj148O7elzCGEXHbuKEH0snm
f80xcG9IlTKWlyepE0AH3CPn+9nD7CmttS6FG8MIK+Y/VKkOJ+9xJ60xHH7oW/dPHXuwxe4gqTi/
Tlq/dQmm72FGVX3KAxsN2CraIzwPIcB+pro0M0hJO0VtIZedacTxIOMDbTBO3ZVXly5+Vlt7ek5F
+NTg6NEm57XW2v7vV3roQnTlLMyoDTANZq4ZD50yiHnfsIGf30FeRHHRSBV0d0P2IThdcuqdTx3J
bsCoZzsJK3KmttUkjlbOllCKXzcfcGNjLYchx5ovwYDhHGDiF2WUcKNPukgXX5XnReygtUie7rQk
533EYXuhc2tzE+Nq37bNuR3VVfaXVqYDLV0fUa55QHpLML8FMs+HYjxGiOb3FlFzMKrJDfiLWJex
HKx6BoBqOBN+AmcljdUjt9w0wW4kIOr5qk9QUtTVmwj2xOVq7xI2EXn/159sA553RZsGSYkJYbEz
dN0Zjc9BaKTBh1GnrWyAInH20J1RyacKboGAbOGHkKVJ2cMYy9iJlxDFzL475fQlhU9NhAQz18Bf
iHLQpywV8Fjt0RC5M+g8pRqi13SWQXsqO4mUP+SVJ9cGoP/R0KbGCJoXkei/X3pDGyRwk3dT0jFs
3FcM22eC570Y8xoX4TjvXx+4Kd9iqlQAbgC8jHX5z6WF9Vi3MSk3Z7AC4canCngKA7E2742gksDx
Tcfjuy4K6W1/o8ZWI7F5qpW+Uu+MnJG5aIibYhIeZCMtqAS2V3kDvUefzZe+sezLZv6ym+iJdGqd
50T3DfezZMngP6ucglg0cJAFv51w+BO6HyX9UhO+a8reigJlGilEfD2J3jP0+1WQo1ik5UDZaj0t
MS4XAQghcAUfHSftI4ikqWLXkEhGO1K0t3kQ0v5kMd8SkAEz95vE9vvoUis5vDDh2ABzItSGMdOV
XG9zbxEc2lzx5QDsuGEiFZ5oEcofkfF3N7pDekAC2Q8jt/yp1MundRzJCHnYt4LVRXsL/jbkO3e6
Sbsyl52TkebnmQkvTOUv/Ip4C3oJG/EmiSGpW7EB9h91MRFLeJC0nijmRZIvEqri2jrUUzN/xBlv
ggCHdgfNd1DueGdW2X6mClFAlYsdwu+inr/6Tyogyq2zrS6WBocH9MLaJCQDt2oZi2H9QUu3J7mv
OhEqfmBRfHCAdevNJyZ0EtxvN/DDbimhWdYYEngJlvYfKThdm/3Rw4dsUAeadZkP6LlrlTnyJXRu
UAhxvhrl0n7+wMKeCG9ueWLh84uiAFhQcFXYTMpdJmEKvceRj5jtlpsEvUqBjlWEk5kt1fbD/MZy
dgWlfp7DBuygBDjdMs1yMJddZeHFwTqxZqTBX0K+VrWoiWkswqsyoAtzJZ2yZ4XjsnKyDmoFvknm
rdM6a/xkkFPFdpLQzmcOvBoX1BZU4wDCP/cQTU6Dm0gYKppCNNPF/9v2IEkwxLV9prk/hjohtV5j
2bdEsgKuREKPaDz+ign/rQMemGRwwm3Aq82kg/x0+8GC0Cb+1fQ/IGdxDA0jee7BWMA8ybKshx0F
4V8ppiYTkoO0phKJSmin/xryiEXzkbgGnO21BvDh+c7MfSh3s3M/boMuGFuV2Kkk23RfKubqwLBw
bD+x75tjOGK2+lb0l/8Pp91TsigAYV+1+xTjg+zI8sT32QWH94pT0bQDbm4/Av2phtRckzkZU2QI
ClrKt/Iq7PamvioKgU6BWvxgJ57KRIVCUNs7QJq+KdA7SfKXWokkmdA8O8x8rTuBT3+dLW4EgXuD
cQspHcfN6QHF6/PH17Uq2Kz+uqsH9+Sa5jlFI7snDW/F5j6d3MT6eU3MAbJLd02SpcosV7gaFtTp
HiBP3gVIfK3vn7DWXHHKPIShjfO4XyZrID9AXmPJzukf4h2ZhruZGeGnbE84vHuZzd/D1BZ+jucy
UBdl7oZE4My6wcojitsmqHy534xaNyvtfdv1VVAEnavXkIwX3QU7uM4tqcKX7Yq120JQmB2AcbZ5
9Nqy8njDS4pM/Sri8rB6evv3q7P/DdADBy4eTCasCTZfF9L8DXoC/0NxBOlQR5xfrAkNZcsi5rbL
dnrvzrE2Bxi84Hgct2L553uZ1YzBuvxiGo3DeeRPZ38vxNzGeE0+u3eQM3wtQ2CcsfTmcTw4WjuI
OYCR/FrJeTWsAlosmKBr0tIOR5bh8rim9Bl9hL5ZYTj38ezyH6nHcLkoHbdEP1GENYB68eX6MDHA
y7rBo1yposqP3CP70l/v9cmQ9vohCvIE/69DEXe/Q2X67oJup2nTnCcbt1VdRNitfLIZBMCXQIiN
iHstZuIrQOzJUgbCP1IhoaA3wf998x1lN5tQudnToldh/A4uV4EOlRdm4U+6EkgBXa5tyTZ6khES
VFtrJuXkPFT2OdSXJrgesw3uvPEIW0NLoVfHX7ZeytthIp3rMiWohiEm9l/c92A6Lg0V5NPRl1bB
yOyi7z6ddrsSpXFX4k9gUNnoSB8cniG9Di3XGxvQPn6fA6gvx5uTWv2boUm03D1IuasfZuEmKnyZ
AO05PgSh3RZVrenKEjIwtQc8mhcIDhA+jdwuCHTbZQL+hkgdw8BiYE5FXpmF83jCsbbnjmnCBsU+
x80ukhGaazezEIdgqQOl6YnbmKZFM+sBq7DZXOBlLJAPWVvd8+HMja9Rbo8Ig7YmwFDiFS0duMlT
qtpHrNYJ4FR/W3Iw4uzTuHQPoFF+dsXALrXOC4IlupICPpGucir77F/CKuuKlTEF2gh7B6EvLteR
BfQA68aixk4rtCL0pNeNiUzv5TeEYOUWjj7IBEztallzspCqMw3CZh+9AYwIlTW40027mc7ujrpb
hDIGcFcKGI4qAshgsuiyxD+kwfW2AYG+K83FlVJoNK6SKCBMkKtAiEHl7do5D6tEW2aSh4CuMYFF
aHgfnap815iTTMYtY68F6DtvVL87Zho1YQYkHPLs5j+omFsfRTHoRMsUCf+uqgDMKCiYNaFj0vXf
oi02VQPL2nYIOph+3iWv69jrwyezvZlMlypFiRgwpR2zR54CLh1oL9UoE+wcQDB8qN8skyEDiMKC
ENLlr6PqpXbCwWWs64s+EgmpMV5F43CYm9KNK2wELHeMW3NVzZv4U9DfEYotE4+3eOXIMYiBDPfp
/jG9z74BXg9B5fFCJGbVZoxEw2muKj/jC+QIWbVis7SdlpTZXnN9eRveyd2WaqcvVbjganlB1wsS
EIs6bmRkyHhkQP4VzWMGbO210SLrtsx8U2tpyVzxE14m8JIlYMrm8EG6nJOgg/VNjG0FgZX2id4d
v5fgM1JbhfE//WHtUCOSlUeuZCKlaO0jZpB0bMhaorAjtgXOZU2c+RbnJvDOZ8F6HlHbs2gSymNg
nbs1F1/Mkdzyle9Rff9N7briJr7NbS26MuqqJG/mL+JzrzqdkJOtvvll5ESVomr7N9ZtXtdjGgQu
h7JMWLViINSUPKJqWkYPV7WDODu/UwRqKRgaUH4KTNx+gLJv8oH8/PFA9We1HtUdxEUrnWtZgzaW
DcRn9BDAjVim7hfOamtVtt8aZNIWMgaMfyKx1EjCJzWR2X+qicAehWYLnxLepTi2PPcMyPx98cLT
votJXepwnwIWlwKCUBt7GrnKEkfd7Osz4F8jpSB2WQLzj73doJ5vK/AdRgWr8lhWuM6Ipkm8qaOW
xkWo0Uc7hkeNlsEvV1yG37qiwc1IhL76gDvsB19fEyaGI83/J/mTHlWRhOnz2y9+ER8133W0SJCL
+3xLJZnNfm9Q8JOBUCNtnk+G45y+Zo7CCeO7rMkP++J8uzRm2pDGBA/LpwNFEE4kZoyy3GQAiK5o
PBmKmkCMDKZpc+WuVE8ga+Fk5GHWXFm7q1JBHTXHm/KjIv7luexnpXXotEG3Q7OvhrUeuaiCbTEB
ZJGvRldSohjigPJWsSFOTskcdUS4BuKYcQQylAtF223XqTt/iyTKLPoRrlRg5Ui24nhgBrkvnJ1s
2tK0/sPwPoVr1dCl2/ysPZwYggHNEtGyI/iYpuzapou471QFsgZCz7E9NuoDJWyp/FC2OekJyR/R
qwEDSAr3ODy9F8w5MDUGaimnXTyAZhq3Lrn3zYKQrE1QG1LuRjOHuGfBJ4vQolWNYiMAo5/6IlC5
bq5kU36Olqhx7zjFLa/TkwGHnZJYBGN94lKgg13h28t9vJLEtffAHWV/2osItLLvu9ziZ8KGHfMd
ca1Bbak2+Czh6Cwhn7h98BX8MGzIvmRUqKk6Z3q24uPuF1gjTzOWdQzY7IjAB0qNw1MlocUcFUuU
NfQC0wct37Befqm5lSVBJQXatjVk3ufbrR5WOIGpfp1L1PJxDDP047VsimuInGNvLhZ5pzYv4rI+
pbiizjlNdGs+6mvmqkEkOqx5EzcK+L/YktJJChFjkL+dRJxPsiEm+3JKu6zXyyKgy9KzAb1XgcDZ
kyZl+WmQyAKTyUp6A4drVbGFduuQvy0T2dFqyxNOciUQKUrRIntOVdKk/C8nqqTUCsN+a3Ozskq/
oxfXK+3NHLD3nQg2G9TFfJ1zhW8NWq9FthmbAl7Mk4N5rmBUR04BI61sshjrkDgR4xuvSBiWn5Xr
J9TznqhtFK10BkS17hlAEwdXBpksYNkfduSCXGAdg1RAulO/CpkOv0dTIpxSw9Ebed4Z+2rFlbf5
MEXoNW/Sdx2Ac+OjGAiTe/JXUSrW56O7zL663q0E1om3jDo1jE/gbRWogGxyUXeK1B+Bm6YeKwqo
f+ixLfzC8ujcaT1gwY6xiNFAB1JMh0VN3DET8aKbDu5vBHcoqHjOsYcVt6F6mGIryt+AUURdK00G
AByOF4W6153KA8q0lWp2xYJ9pMLQpNqPtIYad30aD9C/TThLXljbpf0XdLhHEolLfNhlRW7NRGjj
1LCeZVIqu9Q0ggSHokDIllikUKkZSKhoDE+2fyDC/a1Xh0bytAD3YHTRiefT3M9UTp/Fuu0xWaTR
Me1aE+Mn14APwpeSzu6SVy5vFS5gAs0igtFQh5N/DyIQf+o3kGJZUfaES0SFVSwFpBy1fgB30ofb
S+1Gr4xxtB9BGuJK+jo59fmTDCivFLmNCWEDpzJy3bTkUqz+nL8RSoovzp7E+6GetMuhVzXtqvgu
P1o1fffrZKEgC1BQpyO59HDMoTPHxSXy72okkrXfpIjWc9IoARZbvoVpXHcTaR/gBUQdlPa3cujX
ZmCGTY5crjWijmUdLyskTcizz7+bGTTobB/xRgTmHsppqz/IW3/wBny2bdx4V7eiqbuKdoqeNWbZ
lvjMwBUNmDuzjcj3d3WHFiW9s2106Do2MObqVaEAb8r9+UaLgN9sEKFgkySd6Z8gbkaOC3C39mk0
tePynYC5o1No2x9+e2BI2Ls7dYoIdYthaIFtEN64RYeR1CfV5Z9nEGwxLoqZjgrAnx0n/VCgg9KK
cHbg5wudktDC+COaXkfZX4UzjKMvC0Zo2N8fqX9W4pdynaewq8+A1o57Ec0WSZrae/D8v3ZP+xPv
JtJLH+3mTJj1xjzNLGyN4fYbNMNtfSjDWltH1muO2Ue/wEIAgkVqzitiN0KSOhlzsM1+C2F2iBuZ
bgG3wrBFUD5R8IrChptJHIC6qKEx+x6RbBXAVHodhO4vvTJ7rUzTsU6+KOZk5pHMAPQZgu3VGOSN
s92oOezJbhe8s1dLLjnTfjplMkqa08Vh4Q61sIAjwaSbtbiW59ZMd02I6g1Vox/kRX8+NbpqJEkB
OjB8sBGe8k0/fp34PLextNcstKcT88wOQL5ofzhRzl5+YqGjYQYVM9PR1ZiLMCvMAFvDY3Ws72v0
RKlNMJ8N5t1NDh3qV5zFJeSksd64SzOVPRHEcDMSkEVGmt+4GP3DyYQahq9g5394+qY99Ezu5Ybq
ZzMhfxLX8yKRs7uWezrzukDo3b489WPhhwkESVfDOJd1en7CoQiFctqdWBRlD6x5WXvJsQYsXTlN
dc7G06KgTaeN5S+3rfdSeHbzPEqWOAyDoEU9SUC+C5YcMwMdte4Lvu6k+J7ZtgkQorVC010VSzWm
LVNaw6D+IsQhWSSbGgEwN4zCEtcGFPehVVL0GSr3ol0tsfujok7CoKvUcGTETG7k1jbcWUtQt1c3
Bomy7dWa5ez9GiIzxvkjwwWqIygSGPgMynEX0grKIOPm7stdKEV9T9wIVn5jE8fAFIKUg1kPTJ9z
VBx1VMiTQ2Xq/UAlBQt+vKTAzo29XC+DHPaNq9AYYm9S6WifwwQagkdJgYvSloeg4na3sGCNMRN6
cmyyQmeWtpwh4yuPXrfkk70zwJYrm9Mr3wmZff28CrEG0T425AIkKERRD3XdRMrRBqbj6ksY7MB3
XcRQg7bjN+lAbs2lv8rLWBkfbNZkAq3o0a1hTEjAo0gCCJZIphrFJBXRCugmA2rMuE+JOtUbXxxG
CBFncVQ7gZYYS4JBDxpLxjLYJ98CJsFTgJA0Q1jLXeVNhDwAl7HhS+Ld2HJ6EFBt9O8tM033eL2J
vJbUpm03xrKt7Ui/JHt7yKfDojN9sVHn/5y4fAkm9VD7lWxuuO4KwOR07n22GdID/Y5PokHFkd1i
BCkhp5XI+ARvLjoONJoFpqPbIkd66rb8VnjYwA+xh1Ir1x5ab3jqf2Xu3vUX/xEV0cGQbmiJZPCY
wVRgLJZGkXkYtZi6gZ+pHl8Nyl+yaK6OsCU9/HZsdG9FnA0Ytm2XBFd+3BXgY1uVHWW1PU4SEuhB
hCCVfSgqrKqx8TbjJ8CkmbgL0v9WnKCzSqZr0sVqE4WNPPJirbXMR13WVHiKS7UpnB54uN7rBXSx
RBBOn8lDQV3Z8dwv+abdAjhjWZAA281xbIrcApZMpfsf1Ct+iUBZAfxq5ldR0k/uXgOrIak146YS
nMSVLeCxz8uRYvMaClBdH6smdMUKgSVpCx1iOrObHf9fCJB5pHP0O98D3ldGs9Ji8ULdBWXBxJIj
nVrpl8Q0HclRitqXMd3AZd9zZAfGVbVmV1XeTRCMOO/zltndhFGfmHcnmmflKIzuPTcn54+pkN1F
QvDYCYyqa441MwOnmypsjVFGg2krI4sEwDTvrpHK56t0kl4vJx+c7kbDsaLJR4JzJnxtrTfGyt1k
1b0dPTYJ5XJdE08k95JGfWVhgxRswXyGkwbEeOoPm0lfpGcptakd/mELz/rOkpOof3ICY/P8QTyQ
/TPdpxSNPnQcHEo8SJkXH65lPDkcBpNQY0e1fEplPXW6apXYRo/iQr6n1TUOK8gLN6k+RxEMBUq2
V/c58nBe+/qDz6FYhX0lFhqHJbBG6sxn2BvSut4U6beoUAz1xAT4BzDhiY7208pR28mzZc6ZG1X4
LV9VfNqUI3XzMWKDzAnEJiHUpl+N0nMxd4PDOImHKMirEawSPeVIG93A/UADPP+ngMBZ/tlBqpzc
4amQtde2FuCdNJ0Hyw5gtO/uYfY5YqSmXfZyiwHsTq1rSCdxWawgMeGPz5Jjv6Xth+Q4W/6j73ZJ
eYk3h0gJ1ASY6YNLHw2jss4va+jxEfFKiMKS4Wz019+4KazA+pVdVIAxLmY8Uu1mzlFTZgAib/5V
9cCBNopmhb/KYNukiiVfmCB/ekQD22QkOW8nAFQXcAMpIQYoakZOiUIWVsshjT409mcq2+UbaQc9
/4CgFs8FmqKsTxaBLgd3sUS9KISLSz6y+G58JBdKZgFWCS8ZJxMRl053+GLALaPGtjFm6hPWBxB1
CHXW5FADP48qwVvS/M1JUpkgNh/FcbkH730JHfcgEKQOO4LJMC7tUJTYu0H+kFEbCaGU6wDEM8mA
9XkYkimw/Zu/vYJAdNT75Ca/1sq6gwOQidFAj/vqTzPeTgrCm2zZDpxWNcVDP1XWN99lwUV36kfn
vg0kO9+DK43glPY60hzNST9BpNxMFmn+54JnYEIBLXOSmagz1R8ZiVF/w9DA8hhR2jXsglJF9fU1
/jFsEdjTE68Y89Bu8+4jGIp6HXXOiO9n9On5foxWL/ZcyCtkH1TtHSw1wVgzE12R3mFhS9QxvEqE
IczZfWrEjbsOl7fdLa9lVHR13UCBUD/wKEjOXbw1zB3htNmvSlrnV6Es1GlNIVvQJYugRFvynFd/
blm8e1ku5qdkD1754PgWOhjBegZO4Sg630B78KXCdlt1aOMTPBPi4qM3gWDD4Eic86WSMdaHULq4
S1JNW1PvOvACf0OMQsUdsEiCwoID5jjz839N0ceRqX+165WL+Jahb1IHN6IqdTJm8fZ7Q0r0rNQX
0PBGKLclW/aM/K8k35qM++KrC3Ar8QVna1bQE+OkQ8VmjHnIJ94m0o5y+vmF2vn67d41xYojKHcu
hRdxgWPiCI9Yc5flXFudlOCJ2gU30yY5qpvOdIlsY++OUN1PUCjZLhoyPFNrUDz6tM8otyo64jbl
f9PALzupil2kJMZjdYgXkdvp3F120bAibIYm+0JVbXECH8vlYi8pXwVY7IvHBzlNpprGTXHS8YZp
u+4lL0yB5UfX4qLlQwQvzvctbwSjfiW1MvX6BJwuH4eCLB82qr3uZZVmY32SJ6io5MDUvrISl46d
8KVl/NJygWw7O3/jEQAv8AIYHCtNfbibRoIJZmQZHVmHTu+UliKPlLzVf7EXTK9CLN4UJJvsetg0
ZqF6ih45RNvGOtiyRM84Qr50J6ByL7EeNPJQRk5Ai197GuwldJpEZkCoLRmxIDR9BDg7CpWU6k5d
5U1/XnoLXdjDGhePjgYEuoA0m0+HMJbGZ6l1KvKa1v/Mhifu+fFwJjPfVJKuNJpjDNg6aQ0k0wfz
pL5T3W3L23+89Wddwgkv8iicn88UcJUt0nFgaP/Wgr32eEe36mzeClOBKAibIR2LQBwwEuRxvxDM
aWrIBHhd1B8g2/1ocoFNj8AXA8rGWU6RY2rtuUKIf9p+CBPHomN31qlpVtpGpMXSSURaP2t4A/m6
dudwQ//PdyBtk4lz8YT6cS9CgwcDHdoAoPsfTwap++EXHlWDODCBmeN9PIwSiCcevLkJ9In8II+u
eTerZPbNfbC8jf6O2I4LFhrdDh2wuCh3f3WzD52SCGr2pvfPvgPFtoCV1G2HQ3eefhv7TsB7mLF0
kMXhOergWWNwSaUwqPfEkiFnVJuFWN2+5fgrkxXmxR6JW19r1OZR3/ZhBKjkTstODdpymyrq7OJz
wbkJzkmlMqznkUSDDV77Z8OJ3OdZJKHee/NFGU4hnwf3yblvRRy2tHPNLM+F+5wHj47bUPdFpt6I
HDNEba7J1f0GT2PPImHGY9Py4uoc9F8XbIjO2fBCMHd2HTdG5KKH7AuPopgIci5dAVRX7yTLUAkm
bjN98NAEpwIQIa3WW5xIcfo/+vmUyZXySPEpD7ff/AxZhQ+LT0PHfNYRLiEzAulT3LNOXxnlHn1w
sPqM8/O00WQFzznjWfXfRiNC1R2M94JXuGmDR5m5EMf81XG3XUtXUxkfP4paYNKIzoCQuGOAP5xI
eCSOQW2Vr86xq3tIWbuE+luiDbtRDDYlp5rpsoWqAagjGLxPl3yOJoYRAxw9ysPRMTHiyfgm/sqy
lmRhd3iogBWk9F817kI+ewJ+TEAm7J8KG/mzTzfBe6Fk38ZKDSJNeD4ALd4bqZRo5aZxARkB1TVr
GAyF7xGF97bhaedTpquoC/KZLGg6Z4bIAdJrKzTyKtgKDrYTKt0LMobyhP8Tj4kfIohGSeVYUuam
6cUDZFQ1LgPcTngk1FXS1HPaAEd1+WH/A/HKy+8GuOeVrzL1uP+Ss/L8yr5eIy+6672A5dAKFSed
Xs563yCNEeA0BPr0aXmpDBHW11kNK/ROyiawpi1mBU4UPr1Vkb6AB9PeY4si8RCYIEEXu76FyBfp
9wF8fTzZIy7hKKO5TFg2lfKhqh1nic+3klGr8YjqbW/3UtO1tVPkKwln0SN/kZdaEpBLCcEru9+V
4/gzsndn20/Y6kXE7PYZuWHpRqfcZ7+gTJ6ImjciUqMGnWjF28nhhG5gHrjsF/rOuaQH6X5I2ToJ
U+XBTO+OcXT4bpStUirfqQhc2gFdnC7tXldidl7KOhoyo7kQr3hrj5bv+Uda+R3FXU9LcHn0LPZJ
yhD02ieeuKYHua44vIThX3Mni8S/77Rpdr8//9Kl+MTd3Gvy/B6ZsX/xO+7YXncv2B3vkmRX1VD1
4s/P3uT1omCauMw6vTxGwI05/9lPO7iT0xUCIwAbyW9WoenN7ya0KQEUIrR+yIZFchnpglBeHghb
cAgllridjqgjSq9NZg3G1+IkD+YwJJN1ITXo0l0jOKLbD6zvQotR3GwYN8NmWwmJG4t9w9H7yv41
PXkUS8ydIjACuJFgdoKKbaADs9XYsb6sjo5U0bg3CDQ01IYOVPdOtSAL5tHAl7Z488Kvyr1z1Xor
yVtePKrl9OVFiG/acZmNPzYczdYinGwKygy2Qr1TwY9/FxLrNxPxR/xgwEhxFO2DUS9hCOQLt+C2
Bq542CGFu4LrNq2JhEAl6FTJ1apPdJxH0uBYd48d4qSkI+G3ebvaGpjydvkOqghayvkTxhZeqUY6
kliwAb+f6bwKbgneMuPBZV2dgHp6UGGf5x2YekwTHSRRtlsn+KqcHVbMwdPPows2si6tnh/PXy4F
GxsY3aEppQ8jmDJDsGtIxJ8KEQvhodQRk81N651uTZ/H3k4qKX/Zlghqrs4NAhbhaATwsdfg0h6O
wEDHYJ33m/pjZr/aO66RHubUHK5s0eX2PRd/SOSiPa3U9JoHhKp2rIOZGrelCEMaiy8e1sCrDJLY
Vk0JteqS+MhvZ3uczBmUWPxN9LGckXAE2HGMAoI1UUwITrZyA9PYTX1fVnbNeJxVtUsOpeuqrF4G
91pFCnbiVZKblX56X7r/eNFLIhbZDVdhjlUMqhdZbEYDOY0sNc+QCdky5ZlyjWdp1vVBjFbCb98l
KqfrL1oQ2UTQWJpYyWyjTdhfIgPWH37BjMPmXYDaMKsw6lDZZJMdMe16b8EEN7Avvp//9pIwE4nV
FQ4i004tXikaJf85F8bF/Mbe9+psEdB5lGCiCYsjB2FRKYJ6eQyhgKEx0Hl4V6l0khExQs1IG7M6
W7JBKxK3aV6TU63EYtdaO/xqkgQL4Cggp91+1BsAPE1ifPcDI1HIjlodPhvxDDbxsJUkmcC+D1jb
hU6XMP9nJaLnVEp/28blHhh1PBbQ0Rezt3JLzKHG+ugtYte5pgi6zGbZDC+aShluQeEnVg5VE+LX
loNDxTfmA6455pfDUzH0Cxw2o632Dc8mSnqQJMzkjJE6Yf7Q6QNM+gqtrXKEiH7TUl67Faw0fpSM
VFf1DVSlpmdTC1LJ8VCAv1QXYib6LdeyKaeKtl3GRp79ATFyMX3cf5yGoFGm6mFd6ZS9w/IyrS4E
qCj/Z1D2COSIG81flclBink3gSrl9mbQLAiZtTtUhJwR4Nb1tlY/qIjazf1erUgTj2Y7K4XFdVhp
eXSlhlN3h6ODL+0O2unGXUKscpj+T3ucTLGqmzTFO1qgErsTeTDCYN5lRGA1TgBRu2vHayU6ipJ/
01xT9QNCbis5LqNBYGrODCxB7xk5siwdTVrQ1ciH1oo3shVoOYssh9A48sBCVYJgyAN32qxH7eBX
tcISCqiEJ1T6UQWAo/duKZ5HNnlLTArBw7FFVCJO9Y1BM0FzmfDO0g0W1PWjhbzgIeKAE44t5XRD
aoVi42n+ky+t1bj+0zSqKLFG6twXzNkRDDXZsXFJEidLEU81Gfy2dCwaRnoSAcLSxzdyfzw5zXiM
JYMUwj39fJjE2JZ2rTlZPYNtPhsMl5K/tPo7hiNKdXAB2dgMuqWUCJ9pYyVe6CvirOBVj0/9qL0r
Iipce01Zbr1BGCC05GgsG9nYbnDSDddEJRbywvtYXUxJe1WHbalhmh9THeTulB1XVpl7N6o8f3W0
r+QTJ52aN5iJ35mnj0Dd9w5OilI6OcNcT6y1b3oeUiZQYELBgfbbDonhSpc5Vo2fX6PG+whbaQ3D
PMhhYZNMCARrwUB/BiRiGaDSZHGOnKRAcXWCy3pw+I+JbdYPXLNM+1fDZHxVDJMxqwA9uqtamM9l
1Hbctlni14R9hq08BWOM3IbhR+9jbpiQe6tQLwW6Rv01pRUX4lGKsn0BGel+X1wpOuSjlJe/RlY+
1CoVmJkrI1dyFEmGd6hAXhqT08INUyP6SuP4T6JneCzlZkkKzvIn15GuFuV74KFJxiPYTdrToNk1
h62ZTh2qUs1SsI6BKoGTeoJN1Xvwr/Th8IfFfMEKbP7pzZVXYLumwa/tGGpqLpXlvWRUKVH8yBvm
diw95aw7Nqg7/pnrqENCfbwXxTRimg4bpceyXVkjTKMV0n/QJZITseggHi+5cmJ34CZLpCyo528Q
Qd5mfoj/6lhSq/fUVfasraAA+93VNOKXfVWEvqa9RiY5S+YZIk5X41YoaDYemmXMmoyTZJBRJXGo
t9HyENxf7HNMJ2gQGS6VWIQh4zQyn508vESqfEvRMWYTgRPKzJXVn7YN3llVIEGUcwTuMMNpRz1a
aGoBZppp9TQ+FBI7zHCx1dcKza4RmCL90wAyqSGZFX8yqeu9HMb39cgElNtm1hXZnXAlK85+QLkL
5fBOOLCyXcwRV5m0X2AeCT60ASdSkO2m7hMPClpHrOPJ6+GQ3JK0y2z1kIZWWHgqzWyhDWEX+PSS
+qoXbRDFRhKKytqqxOc48qzkAsFpVBfFP+pT4zTxgPtjzG3P3OX+QgIpOgdKAI+1Bb2e2/00EF+w
maUlN8eZIp1CMhitYCrHbBiPEGGaJ+to/2PFOgRvhPvxFgXwTBl3v19m33vsJwLO/VuaJ2BslUlo
Rnuhybl9uDrCBMPrmsiV1x+v0v1AieKJ0ETFYcIt/vOXOYiXit1P244S9yg9p9ZOIvJa6gKIecwg
vlOlIRk9dkK5ukX1RNYIIN1cUdPv4GqmqRPlAI8dMPX6uGfilevaCfGHYWIMAHsuZ4a9PcKUMhLp
iw2fV4csRGbRh/ukzxryEdQJ1MxuLXwAXOLGFW3tJspzcO5TDWdncD7jcLkhNVMmJkzv+5XEUHQ6
ApwYLIFgP+BfvyJxOwuMCjGXFEQ8PZa8oLGyA3wV+h+JO6fbMQjyhYQxgUtJ8YNj6oToCECsoQ+A
NBYV2wKpziEIEgbc+RTiXW/5GKnANtKHo6XoA76A+9zpei9pPlC0ZqKpA7k2DL6UbSrrgMvlGOZM
YwXFUfvWcKM0I9nbOIdCGydxAlWAjUa3arbAaHY5z7JmvoW20vnSbf4hPEksCEnAw8/JThWm7Nlv
lrOcQ01O2UwgYbhc0hSexSnkko3sXgew8/AFMftLCFBVRo1v38jEgbZvn98SGRS/1gQErK9Mf+sh
iOt+w7CyxYIKao+uBTSTKekuhgByxzZtCLlYv+biGY5iveN+/DVx/h9Mi3Mn/rC5lkKKmsfvBI8M
gYX1KoD+s64ZpqFh/CthqDs1TcjRzEMMYSftpAVS2ltm5Eh8MdGSJJCtt8elSoNPPTGL4v1shVMh
taGts2KlP/71bZkabLPGofFFGMlWu9yD6JdwUbTwYNAofxylkssQgGmyYteXin18hKfZtfJFdxGp
IjWePMR8Qd7aIj8rk6PpnJPDGzS96ARz1oerOn8O2DBZuKyN8xrnsViuP1U7ghvjbVfYdbZ/21Eb
cljAum5GvHCijcJcerzS9DJdvfzpcn8zUZulOmJ06jONdJ/Y9C6GUJ3jVe5DN1j5mZu7ItT0JKHF
xmaa0Ud6n/CnyLC2rUDCLjGAM/KWYLdfVSelJ7AMfItYlrpDjkgM+jW19kUnJRUoS4px7qxhnHgp
Rj1yzgTDWXYHMaEESWdwYQGTF31oATT201nFWy66uixbGiQl1sBfdpEtdgpRjjyOaKj79J63H2Sq
ZMe11eU0ggl8GUr9Nl3/eJUNdkoiWnlQZmGVTWeyLlwJ12ER5VeIum/WBCyM3Ag01fJI2VaipdLi
gwaPq1Wk4E4bacv3B0h5nTzGUiUPn3R0mj6oQTdZrX2eTHrWJu3vmlLt5SnNzcn83j9rA8UpzJWQ
dzAuOE2girK3RsHOoWcBK9BKfqVNwt5r6fWPmj8hzddXanHQu0f1ucsR9Aixt6P8XN5xZvlvZ82Y
p64cZhMDzaJYn/mAN7FJgxBagSOqivhz/jBB33qZlIIXGtNPBVIHNnvm/VG11QDdW/Bpt1jS8dDB
fjIBaOVBTamZW6PM9LwPc6//MxzqfTBnTS/xUGU+YFTo8nVc/mhG27/IUw4437oLNAU9E4HZXbgn
rUkHG2VXCMo3z51t6Wuj6WlEa7AbIJkVKbiLAYYUTISe7gkrs4NwxETUyQV7ND01spgqxpT0yIsw
Gq5j+XZMAge5IltXWVuok/ymOpvq0Au3M9DkgsoRBinHWeNhzgMq9gWgpwiPbiqV1V0DQeHeRBkG
Vkbh3PYJKf01UN4JNLsruNuVBIYlAoxs4shNXgqyBiHI5iFRvQxoRcr3hAjHw8oant+qTb75DaZq
YhesL2usuWf39b9xZiIPYw5Tx3PCmwgGR29JTx+peuAdItulepsOahB8QQk6k1fZF0+OH/3lZ74h
RXUs5H1za9NcH3m+s3uxwUnIcH9d6ATqWYQs85Eoi+7OzVpIoVO8bfCpsnwbA+o2cIdwfuDBmBBe
Ev+MPCrxgWDGGyyDcFW8UUXYreAoypGUB+HrF2vB8jyC167pObFgiP+SEeevgJ3oVZxyzVq4/25Q
G371iYwj43EW7PYPsccGBvZ1qvk8nr4aMeE9KHCedvpvwFpZbKPV9N1g8R7Gpro9gpoIvUZcCfOR
kBmZLWuujJ91UvyM+DUMo9RKAk979C4t9TDILlJmHm6WzhQbylM080cuF0QG8SRqlxP+EHUcvKuw
pdSXcGw2kgUdZEpfH5MRQStvqdJsLc2NBlrK6T8jUU/M+IkxYML/JWA8Tg0OgrLH/P268i2uYTDB
iCs0GhECco8supQ8uuK5T/XrZhSu5NIVLDlweytLSY8koYbbrQu1sHc2HeCHKVuJWYZWcAjNBlk4
eYaYhRtFbrbkADOBzuzr8yqacNFO5aXMNpNCd8X7sRK5uIJCagA1AJDTAcTFwxIcHvWxs8Un5cG0
en1VBdkwL9McSipHVn/8BSpu+9I5lOp/OJFjD4VE05Cm5EVT6rW/crWZo5lQhpbpiHzcJcgs1Njf
n2RVHlCiDuaZ3DODsf1Z4z/Q0RYlBoMg8t9N0AkJHdRHHzphdNfcERmZVu92XQiV29F65G7s3Y+6
4F8MnkLzAnAUuEoTw9NbtrSPw+oFnBmc1CMZzJYS6qQIr+4oaz79+gzsuSvW8hf0fcZD891f7lLj
Icuk+Ksx7p2lHIxzhVG+CHmXOhu3bGRrTo5I7f3N7vmm6Ta3217p9MP9Megw775HvD+OCbE0Y0nD
LsjOuobZ7uG0UEpX/YQFRl9wTW7o0ynq3AHKODEClFZgGgfk1oVoSxe7qchk/tvTRYdTVWK4kBCS
m42ZeXgbY2VXRaup5NynVIXmdqdYrLc3FJjupGexJKfZUDYBMpEZAf3ZsduoSGepBrezq43QU0+1
dDkX8VMBX5ssIqCO9Rord0SOd0zy9RNCiCqTHuwR63TNQuwjS/EQ1PG/e0tOkZViRT8fjJQrZVmu
l15dSnrKtMcBxVXFBknFgqpNdCnzswYoW3AGZeiSPQqu0W5OxGyZS6J/0NhuAH+GMox4J6HhujW3
hKmi1lOr10S1x/cbsDIwexCZy0xwQPFsnFo3sMLE16e7jR3SDgabfyOsDeBq/x1ptcd+XBkhhFXw
sPBmAipYF95LurWcZqkgCZaBK9CUlap8X6j/JwqeAfbzbDmndX6xaXHhCs/vhimrwLQ6DOvuCrmV
irUTgbv0u6EbYPuv5oxYVV2GWde+pts6xJnnAnReSNOHGq38bOL5NgZYC+MC3lVukd1bcRcNLHIi
zM3x9GySdzqR3O/9Wl63/VBdy8cHWX6G6k7gRXapVheUbPpT9XMJ+MovMJSPMhOw859+t2LN1tqR
M2wqEDh5NbVjBPEFGrUjnJSLiiEnL0bRbBlu3ZQYcR3NU/OJN6umg7EL8JConY0J2yxyNp+Hyub6
TJDGQ+MZLS5GdoYCQxcRywygAJP2Kb67H621ITsNfgvTwNGsUIqHpFVH97oqw+Ih75WIXlDhsaDW
BaCl99Z6w60MzEzUWxHeT0CueOpX9vEOEhVHmgxqYh+nxdMZWHl1pKQ8WgQMkjaFe4Q4VxHYziE2
f4yEi86IOkH8G6ILw9sux42NNhDFJB6Hbdw5XhZbvE9Tj9NwK3agVfUQSR6/ecTzbtkyqa/HyJFo
E7kStEEcQbKapJgkHZwJExjSdg6IxgSpvgod4/xLo5goj1FltKP8jIWRX82vFY6FXG7C/J0h4NW6
QjLGCeFkUQnqCvM6voLG942YU0ycRTgCCUR85lOi1jDylVSfF8EpqX/W0wXHma68pV6SSst9P2nv
T5A5Gkecz8Zx+JEqaEnTD4KtB8wtf1A3u9zdxQdDCWaNWTskl0zCBgrouhxqxnQaps+fqTqKRcjg
1jrZPa9dz+RitPY8GBNs4kfsTZzL4Mynkm5E0vWcqg11ZNQfqSljB1xVHC96142CDB882J2l/Wpt
klwQcHzz6v4De1WLHWiyAksdfLccuIJQOgQQZTJig9VUpDK4WSQF90QkgbAcTSbATAcZvoDZWb5Z
380UlFJKARSSuS8Q9eYUimMIjeq0wkNZ1Qmt5ybuyk1bHOHUHZgeB/RTqsbrywOo9+NF3FLsxwUv
UnOw7v0c4KVgQrpJvZnmtttOPaHw+zyxHg0WMNMcOuFEdpG3CZR5Lk6xDs6FgQ3bLuO4MkB9/C3I
3MA9/7SRG6Y6Su1xOPftFSi+UnbTl9zze0wArRKO/KhyGaYnUdgS/PkrvmzT/IwKjS7O/UX1vZ5a
7PUHVpvDQNq+AJeVBZvei4yuxPcRh34oRYRdwDV5yaVMx5h21zKGwvRwNV2aiK4hT1nR/L4LQg0Z
ns/Dn3hP2p1oqbF00LeVmvJowRAjeW8MH0//ecWWrnFgZE5kY7Ms+cZhIaow44ewrOepvRbb1+X4
LOYKFwfkyNizBm48kDQDfbAfbmKJ2GrSIWx7ikWA/Gta8zlpmv05gJ+/pAh++b+p9hIUjCSZOFY0
ZMX5R6k65pdtkKxTskSea4EYopg0k1ZMCBXEhC70hkTVbiS+Kvpk414oNQ+Z2kRYuebC8IefF3vp
a9ge/vMwW2WXO5JXb5YAN/5I79EUyoKc8fZDhqBqrFlwleb8vM9Ekh0rkpcwXsR1x+c8e+6gsXvx
YLExqOcG/YYCs/N+MgC+Ovo3CfOP3hsxAzjJNvGbHaIchogs1JHwME4FFFT4cM8WrrzEvCe4BjRz
kmWqev/MfqM2KHOKr7gUm5CJcoRNAnIvGIViSiPUG4esnSpJsH/cvQQgmRZ17Nr/flFvoR+9bXN5
ETYgZbb183p5jlBm41Dg49Ab6UayKEK/Up5CY+05bOIJwVYcSHeg851h2/aScebkv1R9V8ZMl+bs
wnMm3uo6KjM/dh5wk3Vc3V8MVr0yUICu7Os+gHBZ9Y3SSVtGKH5s01h/ZxOSp7oeG2/mgWcZxSUk
xr49SPrfXQ7oEJPD5xhRBzXwkoji+O5r/UjHoFsjGp8GwWJ4kbfQLkU+EKctamfUNPxK115fw+Ec
TCJ91f14l7V5jPfYgx2Ylcg/w/OLxh2UZ5wFjsJVudMwXcEBlMtu4uNYVTSXIJivAEuOV2/CxBva
UlctJTPjrYN4dUFPFp/Ov4Bu1noCrbvlhyCB3uFC4P9SAYkWkVT1kMzvY0LrcEIewucfedrjIcSV
6PDCzX8l5uwMgHjJQv6XTzfBkzaVkHEYGuQcwQLBsU01NV2wEcjv1DgeQae/KJuQl7opnfaFdZEP
4VbiHieSYPngXoCLYqri0wGJKrZi8UkNEx5dBYymLKmyEryt+0oKt7y6eR57L0TVUTKTMI6QHsb4
aVPIq4fT7MSZlqOVe3efm7ObkCm2zzkePOxIyV5Tckn/OjLVGE0GAKtqZ38o4uUSTaSO9u/sYWEp
f94zVed61A74Z9dvnjwCoK/RXpxieBKXfXscen/2Y2TpV4hRVDYKfU14aykelFuspbLKGDw9rE73
0oBuYZj3vdoJ2pmj39U8P5lyS4hC09MhHht7oz0/CccqW/ocEDtgu9Rz9Q6V+Jv7inQlk0Llge7f
bCBm8n8wd25aF+VPFhAzRNgjJ2azS3fVUAaP62EOGMAevfHJ8NpRac6PfVh8PwCqI2sJKKOAzbQJ
1W/gytMNmkboDD6yEwAz0W0G4XEpDL6vjzvRJo5ZE7W5hT1Bqt81k4JQr1yvrV+Id3wiTnB4fRVG
1F6oKXPxhO49lUkRP1n3lyhQ/XqxQw8aVAykrM2cfAVkvSuHMfcbZ/AOgR6eKpTMfUN+KZT0gscO
p81p1Yp2jd5enO1UOZKqFkQEqJmnbsaAR2Z4lSE9vkMEvRASgUwdfFUVRf463tq8W3pD6T7ei/Fz
jqinMLyReczyMHtZB75FReX5TIdh3e0nG+OQg3eFVomYI7VlVHw5DmBBIthLVPbmEdDW8jWYutY0
4zhOIPQnUm5hxHRWWTZbe8THgJ6YWdPHSzFP2V9vWXjkCVDn27HIflKwIBLLCSVyLsUap0jnLjbW
SHNdRXzD0dH1RdDuABXKLjKoVQQrFlz7u/F0pRL8HPUa8DLr+dQnxQ4AyWob65Xk7H/vJqxIolRJ
y5A7ARjnC1Pt1vW0KTpplkOaw4RJBl8WBLA+w1D9L5DzYo892FLFyWCt7aH+pC7UzjOUWvCK660I
bLd7LLNDsUjBxw2+Jd9kNXsrifCIQo+jX/ZKFW4PJMxplSt/IHVZQfAj3DUwQctbXKcXLWPs1aGN
mcwVIFdQ4unXGQ4zy7PvGNCdMxkRDVCnVNatCbhOLQLcYw7dd11KgMSeaSWIu6yvqzNBAxoM4GGF
8J7tidKEgV061Oi8JPqe6DYhZIOI30PFh58f6v24mwaK5tjoIueDkV+86Xj6MgM/jWBLXc6zWgrQ
A8eRJkW4QVWm3ABWw/qB90hOHnSQgZ6Yl4/Rxmuu1uIiwpyQpmy0hxR6pz5SJAQYusDAVQuvRNPs
MTxUVfjZY9tWAi7yJs3KMwEaZIgnbgCHjBhk05asZ1I5chVeOm23FT4XYmeWjiTYSVTka2mtXOWl
nVoeu8c2zludkCkJqjBpSSZ8LZpo/ZSAL17+SyuarSFyqU2Q3j9k6eD1QJRLYpLh/Wb6GvR0WTXm
sZhd9jx2MNl5wcoF7iYLu/5vpPrQjOZSCine2Y/HrOm4wEExBfDUfviesLQF5t45ew/IpXEg6CwC
BGXpKLjWacxU5YLxCOpjMH6LVw8e+6C/Q6kxvENBev4IgUZ07RDCFA2sY9SL/NcxcHPxFUmfPuxs
OoKv8FMsA1Uy9ui7Jw2HY3fWe3KPoxMMD4XVPNz9iUHkfTujAsxv/kS3x4h5mzsQS4vo9Dz+Syw6
w5obag39FS1jf8ABdYY8EpEfvQhNOQz2t4Zb5iurTrKEFKRI0VN3Sa6Hwj7RsD+zSHrwl7W//xqf
TeUidBYmKhkiJGWTcfzc+s5flvCuRn+I64UBOmM+7choGQtK0h2vKOk9ZiR7uy1FXHDQPBHLBf1E
3eD/rt2Sdx+htIeM2XZcqllXL6pWa2siUeOQfG41ng8D28v3AHaruTxA9rr34QjeXwFgIk27GD/5
epf1zEEs852v0EzE2VhLyIMnaoZhr4cDgP15F3OzNBDJQAX60CTBlnZjC3eABgPmsS0d5FhWz2te
uinhv/gpMMdMNLPtwdbwvGXZS/E+GmyXwKgX28JSJCYpkr5numStwaP+WcAWxQEcqFpuyLLSWfHr
ZrPrfjLrra8w4B4IJja6WRZTaeBuXsnec9fDs2lcgcZ8oaSzrLWi0nKZ83LNoCfIHIpsKkt5voKg
Dw0NEGBFnguMLbaJdp/WOhBLhcHmnTsfozNaDYPCnMJn6NV+ffpEAklDYzy2cM2jeFn9P3W/Gn+q
F0I+Bt+WTOB5Cq0MwzfwGY+o1sDQPmKX4dgOmTxz5Mpz1xuoS5TbAkOa9t+8SmMTwDthDYrEfjQ5
7GdwkghKjyiU8V/crLROZSHcKc5G0urOetFLyKRh1Qc9qvn+czpyItKDTWuY9pr9KH3e1YqgCPDJ
IjejZhqhd6TgUCmeoMhdXEehm1i3rMIThMtslOB8KMZtuVVNdyxmeLat3ugVOJBQDkBIk0pb4T28
9K49LSEs2DS2bpG2hFwyyK3bzOHe3Y9mI8SCceBwfYY6tr4nmNie4fXMa6uJCZC0X7sB3qki9gma
PmEphEvBbKbWjYamOaM+7a7iQrzfnRy6hqvlGe6JMy5kKUzE2LZQsR42b+FZSUr51Vr+bdCyKbhW
o5GrXOaHIoElK59gAx72+REpBaxRvr0fzmp0q5yI16k+hbnNwn6EnaDLemLYn6/IL40roI81jjcO
XXqoGpPZoA1mmOiAJcW1L9vVf4XRagG81xh/nAm1z7Bb3pCSXUqBNLMzU3wWQ/tr1Ts5VYZpS9e+
sjNS21/ejMm/Ubu9uV0zd5fPhtJfeVUlAC0TIMapP/u6CROPADEXqiAVutvMz74pcAqc3OV7dq+N
1KOaYPV6LFTVDNckJjgqPVLJowRTnlvBF8qZAB6NL/egSjOF6GN3ValKKVAhl/ToRqJCeXpiGN5V
VkpuBTLel1+dRNABOc105ZQgj7nwESFL+d/nYpy4BAhV/52lYEC2ccHe7CPX3DUWqxmLL6JwgI40
SchFDv3cr7V9yQ/0DC3/WRfuz0C9p357hq4mxY1MNc5XPB+t/gs6LFLGWUDKGl5FWcU3+MbChFuU
jVRd//hrn7zzQBpqwgCVgBS3CxayeIqGPsL/ia5Hp91Q8ur4b4zBsoL/VdGU8IRVO84xDOzNFRSD
RL+qSuqzeaTyQyQo9s1HkxqB7NHXe0lpiLvNzRTQnnNfSVeRDnMBPzMqo8d7ud0ehcxzULShxgtf
eZQZnk3oQ0guRTw376yb6Hz78LVRpemkCb+BDmeJvNtwWoZKyID7wDiGb7nlRfGrVXHBxg/9EGyq
5WXjep7sJow+lRAXdAcnKfp5vH3MD6BY4EleUWktQl2Bzy5qTxp7l4JF+ppZGgozNee9QwAvbLBj
Pg+xYSEHdQl4u3GdfOkRj0xYSe/u1Tz7ot+2JfUiHrWaepgdr3KZZktjoK7s7dXY1ZtUPDCs8F0V
VpBP1L5X1sSdGLSlnEVyc7hg0iD+JqZff3qGoj6frE1cyGRG3WvjmAvC4MrbTwT1qcfM9BF75LTq
a8Y+tVV7DaS7zrraaklsVTZObdEr1HDNo+MsugAKmPVTdtNMGuPyELyl4xRDpofSy5Yu0YjnciBD
Pd0Pn8FHnsRsK+REnJcvwzlu6t3FZHmGQGdSid+oNU5Je+rpZLSyvo5O9Rc89nMHI/6SmtrU1gc+
TK+xLEpekQWvaHg0cg6K+rMWC21XIRu3oIceq3OfcC7leUqDWbE4XdJ47wQICNCRxYaFHxZlscEa
AxxMtRARHu1y9RQ40sxyhkpMzs+mTkllhAL76WRJC5w76SOBKnHe2kz8Jsvwp/qwYNrcAeTXVpFT
Yn3phKNfJ7GS5VnmX0/kiDMH8SI1KBbRfQru6kJo7Z+Bj/ILsAQHIZaz9IQvOxsydrRphg9RLVpe
3nhbnD7c+xSiLDzEV3eGKAo2qJQvel3EFyV00oMoQ+4b4BzhuZH8Y1Uq6tdwoQbLsvxrFvN2QT8K
bOKqIrdBxzeqTyTYUnFwYwuXF3gTcvH2TkDNpNnCosOJUtR+ftjmznQ17XdexOs2fy7+C/4Yy374
bIJpglupOj6i9yhD5LaXvNZNvBZaAI+hlebhBPRMIiCfnbw+zyKToO2dIx6bknd4/X3Vp8Ykra6K
K7XDYh8Z+eunlMXrZF/Do50xz5uQ5QmvWrcIMu9Cu9oel1spSDAUcWfYMoR5dmj9oLgQmzYwJBUy
K7jsBjQmGPn+uaA4K7GZS1x/q7dIRb+iVvt5iC9YSRc7menLnIhCcbEWvYZ90dGytDvkhNRoQxZv
YZbgajnkKQjIFNJSEMVpLIH7gbneEAiRhITFt+QB1UxYt1XLQ/EYQqzCMuf4Ozgovtku+DhaKkDU
FSARoFUzrSscHWQEpn9T3JFG/SZOq73aQ6i/cUGtyt/czryRbPtR6D6A8+SQ5t+H0B4RpiEohdbj
NBsCrH7EZFpk5HkbAngVczMtooogaQRSWqhhOEq2gqXn2zkwKse9y+vuvIi7SiL2lw08VWb9x4X1
bj0gsD7a7l0HAxYktAQXu4JsAuDBYpJOJ22z6cfb6dpJWZusE4jhB4W5xrZdVmYJeZCZzOvNju8x
2WJGTmoHpLvnK9Sn13bvGyGeS8SjvPPiP7o6SzCg50lZWsi49b9KxC8ccY5DoGFdmlcJp2a+EWsX
w9aN5TJTlqGdkDmMbu6v56Xz/TqI4sGjvYuS/pJ5bJB+lnM4OA3bfOgGbNOPcEc2ZncVF8/jVhrV
yqMhmia+DDkZOgyUu+KVH2paLrGXBNE3Yw7PFh8Pb+byiG0HoUN4Ad/YaQCwZrAphxMJsWI+b6Om
sI3VsMs0dZ/IN6Of7JKeBCrSiLUkVLJXm0/LMEnFBxepFSfM+rEwWQ2A9BJGdhTnoKqmUNsM0nr2
sumQdXfl9LXEio3VBs3xhcEKZ0sdQc7beFY0+p7V+ZpfBXsDQfc8d08GK0c8+XLIBxS2YhWkq+Bf
RsEeSCwA9y0OmFQnLhfX2SkkSg7M3LF34Zq63BVIxrET9p83Ngp3L5ufFaR4DwBhYhMenZbUnpcS
Mpv0EMltiT2ZkjRNne5B9EA6EBwWT1jdgY2j74unQqwCnSPjPu4ftpFh/7vlFbC9xWJjWpO6pb3h
LJ3ur+xpBYatgp28NlWUGr5r6howVXjYTOeVG8wmHBra3kIu+mdHFGFPVT5Ohry6MuGHNgHoQY+D
fk+SDgHDI6KeuLxAyIpxcN1W8FxZP/kkP/Aj6AxF7GqUtr8hfzkPRvJKnUbHcvoyNN+QLNJs2Cut
0+LrfIsyZcj21WE+A0IcRAi1afeCr2sdeeHMFP76eQ0BsV0/r3CgZ+8XFq7Dkrjcfu/o3LO5bBUc
W+1GjSDo5/jStMZLn+uRBEoxKsx4nDNh9QBW7Cg1BBKT2ouijPpgFptTSsSNhtx0CZHkZl56t+3V
Dd+X0KNUbxJ2TcgvILfgRyYaLQt/oALQunAHALqzb61fm2i+KDwjCNrKs6w0sYiZMEmoWErlf63u
4gydS9TEWR/9BYBiznGPEISzsCyIaDW8XlcoYcKZ9Tes8Lxa47CFrfuYnWph9vqEWlFJS2bJjIv9
Lu2en0RQ32jnOekOnFwD5BwXQr1ve+kHVKdtATcFwkND5Vgn75oLTmYbST1JGgw5k2v3085jMmBv
3kDND2OysnvwV/u1Jfq3BFkhBjWzeyymA6CL0Q1BPiF6rItiyv1lkw5VimFBtMb/aGbqKgGxmkH+
YUBNnaIePpW+wdR79+YzQlne7VvRoPURzb5n+7EaIhD5Dvg0ro2IBvOKIhmvrjC2yX8JKga/WGw6
jTwtRm6Onbjz1fXl4QmhAIttYJeT0juvF7wMQq2Kj9wv+g2ul0cdGOm3OafNQ1/fsi/hBjcaj+ZY
CjJCTxgJ1kslXwlS7PZb0VtyZTtXQo+beoz7OTgKXJAtvvABsCaBFDmiEoOKaHTh9hBF5ElpWDfa
CoZLbfYhU/zzYn/go/Ohq38e+Wrgxe5rYV9QKQdeP8E6dtijOdmE0KJm4qfvlzXNcnjMpOf94icp
kthNoHod79hVgP/0K8FBliRGUt4n6XwJXHlwTVwMv5aZL/EY50iHm/Fe8wjYtAohiHorcaHLCg4j
bwu7ZNKr7wsYPCqLZf4skwgy2pnSSuO8n/VXT3C4AljbvONwkF4Ue1/x0OVYcRfuPmc4++SxS8wA
+cfEr0Ehr1BuEgPbD7c9+7bLmBL5yTNJQ2qNRSY8KOATqD82pFgRpJgeB5OZ9Vli+Wzzag3y7xYo
qVASgeGaiUVKPiigIwhFO+q8oBFwVr/04EeuZRt+S4eFwe3JGC0Q2h2Vb02VR4C4kVAuNYinCxxm
xnU3b3zZF721ziH0ZTmiLHv1jDSZdfXcq1+qehbP8b59abK6luQ9gCCBBoiJfpplghYjPOp0LqsR
5GtRz3F0JWr5JEK0GMOY5Dloq5Qtiq41sDdgFs5ntN69tnzClXnYAbJcfHvZxiC/8fxT3+XHE1U7
HKXUUdVYKp/elfbnimdn8N1o6B6JeaGyblian9i/WzTH0ktvi6IItthVpnnidBDFVYWVHqYkh5hi
8Uy9qB86uyRBYo2QUjactbfE5SjCS9uhBeXlnus33vech9LT4ynpoesQb2jDLit9bxOwPtW6l8fb
Vb6N5KJYZKm/Y6iQnRE8Iv2102PTeqAds3hyaF+yCxAist9R54fIb1ri/vg0IJT3gC4rdWPY3WLb
Rf9PP+EAChkmMxX9tPFM62dndJvMScPR51bv7VF7VXgTweNCKED6hzPv7xdjxgrAjB4Td3+w/bWl
dbUNZMzNYmFXyxtw7yOMouFh/Y8HWcCj3pc+wTuGaEPpZvl66X9RgQ+JGKdxXhbCL5P+t6o5Jkmr
lZbRI7TgUPvDntNdnbvokdl3Ko87vq8qAD1IM+DpW6NbeztFmP2AwlnzGrwwlDey68bAO856/GgB
lqEOjbiFjNYQUHKYCeCk/IHtPVsKRpRd7A2WOtQw4uJu4jr4btVavapYK0B9XZl/ukXKUmuJZu41
j08rvZ/eDJNoNvyvag/f9sQKiNtXCQ0y5/ekt/Lcf6EjzEKFo7d8qbkwb4ZT+yrsactQlB0c0Ioo
YkT1MchsOBNm4xBspD7JuRtOOJy4DcZsXPC2qTAF1M2MXoxznsL3JnhmOE8ot0K6H2mDo/8vRfI4
Hz2dorGExbNi1alkcmtQJkBMtKzUByXPWCyubWtvTM1DydzgSbAfjdO07BXjXAgsu/+3VLdg+x1n
vWE7Zlx9UmxSOcTzs5SdvHbeP45Y39F8t3Bio8O/Vx7MqSKnqAihEiilko8eU1sCmx/ybPEOMgem
rVQ1PGL8lwvJZvnyd/utzzASDTWoYyBDaXrzFuVSlYgPfCJmyVNxxUkovT+ruAs0q+Dt4EFMwMV3
TZSZYDk5K73aRgD2aPZiUkY8i6GH6fbLE/4oDcJOk4tXBVBYExFKf4PloTklePfHTb7sEFnfpC6U
3L4bikxxkt8+0hh6if5J1aN0FqLBJua4hNgBd3rPXYmWn3E/IIBnJlB6vPCFAOkrjKPTdLmT+8nj
1bzoc703TyF5kUrAUhYbAIRYEZWF9C227miFhCYNO3dFxUWchTGAP6NaC1R7zb9RM/UPEYrpf1cz
cXnZ8n+R9h9/epYLcTKB6ui14+IqK8ZhleH2FmZRwjE3a6cDL9oOzJQ0RdX9cIa1fiOgaL0CeS0U
qeVg2ol5hnfsRs+6j/d5KuIzMc6Ggew9WuE3lOyH9q9/b2VgfjlSKgpB8hMr1+LInXcr4nKzpiEe
s4YaZjvS0Cih+V8wL8Ch0ojNWz1CaoSx+mNBIuXOhzxLQ4h9hw8sqxEKhAowWUG4Ki/FqSUFjGyr
/YUKmmNBDPnktV9oL89GOKVxjIIlzSeCwxYKgHRBgp97/N5eSKX2ijd40iR7zKxuYYOs6iIFVinN
xmdt1EStQZv0BIikXdDQRp/f+bzecKYl07bFiGv6SCK6U0WqEffigeORksphrSO8FT4gT+ySuQ1w
6uEUB4kqx/OXBDnLbZJpEUrLe1fUUPQyo5juMxz49pxb7t64pnbPop4arJBEAeCTMAOCm4iTycd1
wipQo9G0Hl8DfDwbgsxpba2JgiYUR1Jdqg7D6RM95XwYXhv4QhinbSlcSPUky0NQzkxyeE3tNhKQ
f4Z9yQtVJ0VV3EG08yrfqZw3R4rr+pbIyfMKO6NBWaA2RGilKIE9/eIuEVaizW6IHxuOgp6nfi2r
qEQbVbIVttPV2i54N0hf40VHggVkt5sdYAzqa6gCtPdXmwOOGfU+ecBKyoq8qKG0ioi/9053GJDo
sdgJWLnrtfeT3nhYvNAflwzPO0euRGeDX+jd3EfjZhIi2XYy+6UzbHgj80fU40WmW8NLecAr7noG
IyEZ/Bgbbs0XuSBmhB9AXXXVV3PZrEBQVY8ugLIT210K+ihT5Ww9qaJn0Z3E3ShZveygJBU6XN1Z
Eqlgs/leFNldZvK9bbjSe0qThHo0zuSadE0700Z+I4fixgTH1GQBTU81k0cDy3yUMJvUyyviRA6d
u4M3ZWqtyL7evo86b0S7CK0e37bxl8gETHULwHxZLeFqZNvsReguNnT3SrJqAXpx9XL06b6m713l
yuKfT6ssyMPhkJuZz6ksDVIERvt9/osfsHsPzJF0rj24Y4LolEX9RTRqmrqR+vh+5N/8C0uZnSvr
3cllTXvp3BeyAf93y5VHtk4pGYarW2FTRW+pCyRfbWq/6AeLraN97qxktuumkUxvGqkXQFSVM/Qx
RsoN8cfp5p8MxgMAnNpuscQLiQqLrd7Q3yEIsj5hja8FVHrRAlqNR+i1TkGbQDsJv9+6WzIVY5Vt
3Xdr9luhNSnaVpcNIcsufHgVo4nvwUncQBEvrlSc3uqhz6fI5TsvGzWfTU9uPkohldIoj7Xmvc6x
LGmrP28sE4RrW2WOqyNbaBSy+++HbG7id4h099otqe8hOUS+BwLy2WyTJDZqmpGgnRSilKV/yHP7
wbFTO+1w6p74FjITXLhAqEqlwGJ2CPMUR+6qDqHIdKSU6dUf5XSe9Oqw1Ytw8pJ/7H4C/NF6Q8Q/
9ndMh5E3pVeQePJsZhcNpsBzLzEgeFHQZOIotJKgAg/YyqxW2zkLhb9D1zz1hv3WA4BwRY4dI0U+
81NI6+2bDr4H0yJXznHFrjRvizQiVkMOab98oKryoyqut7u88Mti6oDw2VyMQtYcOiCQo+zvkHNU
RTsT+ZngOpCORNv/WsSRxwSs4bE3pCwY31J37me9fmCxBSx/kYUy7x97vonfIFonxrByl6kBXR5c
hb8CpGchfJ2No0fJXaZ6EOi9Z1mUi5eCAvKj1rGUYK3Ci1Gq0z8AL76cWlMKIvZFxPMTtb5z6j2/
EpQJmF73nkSMKF3GJSjIRWlV/RWRpIKV22/rWgYS30khpUrv49/K3iHw6UP9xMNBEAAq9lEM3ZJI
m6kSDZtKf5xKaBdbFPFCtendBYy7Sadn1MoD/M6jbheX445CMXGk0GuOl+HEn1CvEjkAfHf1q8pp
vTFW8h93Giu8/5sZWlVIig4i87EzpFxTMMO2gWYCTXXjvY6ud27K0Mc0YlgBcUZaqxf4tvPgAOnf
cyQ30FabQUAoGAYZ+FnnnjOVdYb+icSV7vnZmtVibkQ8xUVLNJzs53HDPMuYGwPxnzbdf64fCfHg
Zpz1sp4ffR+h5YHQinugPUOUzlCMEK2J8e1QYnGUsGgnpPAphOPj7yY86kBQvcnx62ZCv0P4BerJ
AbK62VUXG/53ujeTOkqvfyfpVxYBwPlGgZOwLo7B1Fdxl5gbKJBwq87xAUNnZyerIyE0lVtTYWK8
510UtVLCAH2ylj8OxT3vuxXngFsucTDutw+3j3K55yBn06+q4aD5+AzPVRzSJ8B1kyElDvAKL57K
5GWm5KDKc0zt1N0D1VoKAGD0UfbVahP2Yt67jvFTN2CGwQ2Kpt6jZFjWcp9nSHvgQFfHHVBhA7g+
6NJ1yNPWVAS2dShmPdRRtJR66KQRQPwta66sKz/mdEB5CFR1DwAsPfFrltvx8zmAq3UDYmqItLTN
hpDAbuV0yXHuASed3F6zJDu+XVm0twYsoHFNOvyYMRUKuoTnnawsxAP2pdfuap8p7bKJgLae0rBb
1X8v1N2Uw4jFz/dzSifS9xBrrgm0N0KHZbOJWLtMQGBORRSohxtFsXdlJT1DTUwRhHQzI6n/Ppya
mVEvNt2FRu0dszPzrvEgTYXAVU1FRaIJq46NHHgScTcvMkvhW+EGm714DtEZwJJCxZLjD1KWj2oW
EG0HTyPFFckfBa1Dbu9YlKD28oMjOJEZ9X6n4v/mEIWyO2m8UN/rdKZPNGPvn1uH7ci9zphhdWNt
oCqib+lGUpAWXrAkw5IJSZpyNwn3Tn1N2SAMS+y1O181bSfYqulUCVaIeSQ8YCTpHaBsJnXNO7LB
bS+YkkRG0RNSCbP5vshPsn52M8tE1wiN3QuvtUp0gpxqfkAyk/vEEW21QVdhm/Um920ZBBlvwgQd
Iweq5F+UP/X477TRm2jcmLOD0n0xptxEpoS6V8O1lD+Jz112m30PGmBQ5bri6iFa7gEUwlpQQz79
mwlc/xTo41nj/gsvcnCnThu7tcFWB28wfinJK7+Lv+ZnMslTkpJxkw53f6TdKfbm50OiiZE8OTv3
Us94BZfZ3M2oyp8/rNb02td+kRCjKaCmbm3wzo9WzLkWYS3kca5Q8d/z5OXgMPCmNCFds0b57K2y
LXrQpimrd/4YeO414qiBdVsQCKwjCpE6QjwR3iRC1M83u0ZCql/56MwbUZkAGYmELzdgkjF5ZNFE
OSu/uWbAdp4dQnDzbLtvRhBPkDbN67dNFx58+MajOs9CbECYIcV1oGlUCwiuz4c6GrhG10aIy38U
jinFF7MCxnUo0O/B1QBPZhk9XYX6qNgN5MUMCB6Z36G3XH+miDBBTdoq2B5oZeRxMsO3DAcoIJ5D
xOdL+xcuVFK+5iacdYX3zi+DDBoavVqp67L7cid+zCSvxWq1CHxliH6sqsjiumgetQmfMtpSes9P
Rg+R2rJB02Lwjd3SCkT7NYerfhQWjqwu2xZd5lHCE51gipIKf6MOA4HZGx8XfDD7Of0/Ttwcsok4
izf2rN/4ZH2HdM6E+0MJXzVYZ/hVYb1MLaJS03H85CP+iAmBekKX6q2GGWc7+x3ggIj+ZdKUGAVs
r1hndn/7KsxWmaVSgytoYQlGd+io5bBCLFrKfZTHE2h1zzHsJ6QWghDpW0dFVHg1Wu15ynuxcrGZ
9KA1RB+gcl5BcxntJFTbHT/xYq+Kx4TMYQPBVVlS4wtr5jIuv4fy46cSDadjDVJ95asXXolMJJYc
6mHjWIbolvvnTn7ls3ts5p9WqbLWu09I1z24/8n4wFnI+kkaR/PjnAfyvOR+BG0NDVtPaTyf4TNP
C14Pc80eRJuqEU5pJLYr5pc2ZrYgixm+w6bzn3cdJqhJI5keSA8hoeMRUc6biCzvjgksEhvda2lh
5hQlKGveFz6xvdgqziHvRcNJJPWCyZ7MnrME2+tiJ4GpF4Y3705PNpPSkTxTUZfACBV6W836RF0e
crehHs7Ul5RwQAx3ZrWFzezFjVgdUX9u1EIGx3u/Ygrb3ZuUCTPCw8Pth8W33GFq9iTAfzRpRfGz
YzU6yw0sFgiZ0BOXcfFNxek02Mr6b7lWN5OXWwjDp1f7apoKNjK2C1ahKbU2r2WiepnYSONRdz6N
j78CiYargEFKWTGvzLk3BAh2auc4unbmaVXEtzLlKpZEYkvm8oVuhaRtX9KfZKUB7dcV67C24YOH
owoc4L67+/sIhkdI6+Lsi4ENRPymbiXN5fYmTQKaBkrBIBF7cM+Mf7VF3mximNT0DKQ2MhSjBt2o
iPQ13Pw/TOD/TXwBeDcnrYWpJpmPq3yongCWDf2gTWPpBv0vBNaAePlH9vhku8aa3U8dUyTgASSt
8ziYrmkx18XwW1NqmeriVVfLBVSX+xyXemnt0fckDyBKLFZhf374/lACi57C72gdTEJQSOZdXtcS
FHKv4msitd12IvSVafyw+kxU8SD6UcoHu5hD3RTyJYpQxuVYOar1W+HMPxVIoFqpgUHo+mpqZhRH
J34cy2z2OAe72TijGIjWi3xBpFOwGTD5nLlGIO04ljoMstriKxQ08JVgLttzIq6aW+n1vMh1omCv
BZ6Q09ZUD/mjmgWA+gYsYRUTnCaHOmO0ouoxLPlpFskcLP8RRO7LXeG12qXYYegDdbMEdukWFcdx
J29/X+S6fmZhPCh/b6YfqdxoSGeFGbBzc3nOjS4tktxKbX1vNbrSofLFrf2bzGaTm80po9ngTumi
wYX671mvBP6hfV86JqvMGR4pbXVbsnVFFzHlQG79UKoIbe2B7aZWcPS6rkEpC/dqZnSRz/I1mGwu
zwugNT6j4GfyDpeqnTrrlm5yNsnmQTE1n0qWBFsN5MboxSdUrmq7Lrzg14oiTVxw4XFoNZgNeehb
ZkNEQgTUdR64aLUF2PcQ5K1Jk0nGx2te+yX+EsySMevu5VDW2NiBzCxADVW1K/SXcBeu4gOzbJzo
9ep3aCsRYUJLApShXo1HVbzwOJfGlWqwxsbIdnphQbxYVQXMz5heiQeX/EXSJJxX9x+tOuDYnVTR
TqIXrIfNqrNSQiA5sV7iQcaSsfkYWjbj4aO2uS4qKTArUkth/GTgYfrARfu7eY8nPGQ83hV25zku
u5VRw/Jb+HaKpgMRbmHoqEqthXl6N/OUVIiZErG1qYGyoSAQ2wIprPKeaVI4S0unol+ccpIKzedw
vkuiBwTjf+5tE3dXPZ2nD9KPUiBwIvL/pyB4VoRRpQ/LZzPVHStDKsmLkOpoEtDiwKY/MQEZxpr5
Mvg7vap9GhtvUeJzgUCpYDmYPAk3UrYrkYgHUvHVVf8BmI+FBbhVFXy49LwT2OA4MrgIrZ53euAg
HlpOv73Pp9AWpDkSA5GjKqslzgS2A0zKIMxTj9WBi8jHcjxzqezbq1LFfDf3As4Z+l8wewntB0rc
WwQLmfG/AsAh17LcPJ5Emm+9KtyjnQDMvuTUBY9KkZa5sadgCWOOdlWe5xqBH2i7thB/n/imWjGF
LyxHTSi5keh7084pzUGGo0/PaM+aFtwhLk7KbDG/H60cc+GwjYvD50qr/uN3wfYpNNzBUNxseSnF
BDDl+R7Kioy0PLHTuoFjSd5ie5yDB+IiwfD6OMHrRjQn8E8EdIQWEH4OzSX3nO+5E5a4xf0qiYa8
SH57bDVSKVIOY+cpEIFDBgwce4hM7xxLNktX3sI9K2wpFEmdqSKEpqub9CmZzUxHy9nYbqNL/NeQ
f/GRznZ4g5d2yWnVLdsSVnqaNieROgs9G+aobtYMWBwrWaRvxk7HAt2qwvyCuTy4+VnKRKu/vjn6
ZAY0mGsdLQ9lDoImBTW43LGFzV13n5RrwOdWH6J3qFf1ch/6Fc/vKQBd5fPynUoTOjRyukUB1hjf
UcaGgm/FSSDqfSYtdLQxVrhTcoqJrQMAXkBl4KnrhJqioqHwJNtt/3YoXG8oku4wM5HU+bD/UihN
jT70ALvh1C9/Pr54+gJ5ujbVF4xk9yuFRLj4meZ9sOhyXdBXl1TmnPMxjCjLau8yX0b1TjsuSmN6
o2TWPi2bg0bOMLo4O9qs8yyU6bgZycL4nh5RWVxPs+AO07q/vncUUzqvTZvnGSlTI6KixdO7vIri
Xw/ZTm0eszcalXtq80BzNnVLx1CB9xo/++lu5oL14YMQVBLWpE3+m+6aph6rcTw8tsmcOx8TTJMx
rAwzOHhouTs3QvMrgalA2dJ302bFNMNpcxDmu5hUQHZpJpVJhoFd3OwGld5ZAai7YAQAiVGd2Ggp
p0f8PEqO+7s/WxflHEVB1IXtmcrw1I+XGujuaZS1tD0qYp9ywSjpHTSvM5UhhrMC0FAYHEQcohVA
bCJK4lbSztanvozifAnyiLO0RwRT8rPo7j7+/2O9/md5Ogv/XXYyibfiUpZcATg7IlsP7oxvQO8H
wFsnZWQ0V/J9CM2/na/9/qrJxgOjjDnoL2c7dCYOaJb/4WMNgukl/4pPM6xUWBzK5XiN7ucRNiGZ
iavT4DmOWDk4HIzF78x0hmaPpZ9dINcBoW3uiGnaEfZO6wEjxXlhARv32H4jU8O2DY3VGhT5azmx
b1sRkKefydiIKKWCgc0JsjQQcvKAwUnHnkqVKWWRu0MxjX4Fip4ndJOaD6sVDVB7T32BXepXpoCg
iNUeElvtZjwCRVN/RRpd3bcEvxUikLI3T232XAq9+1d2bwpp4g5tfbr1540CXeSHi1AlhXse1J+O
PSGyEELi/bTJ/2BD731J8DC6R0KscUAKrWJdCOcTP+txU2OHiL20rSQVTMIjLcuylHHQ1z6E56UY
Iuq6hEkoAqTEDTSkRk9ie8j7PJrswaK5Mva7ecNh0+vDBEE1ZWDfbG4IkPm2QOEDpe4lqKEEua/3
jV0Ot3yi63oynXpg82Ov7Pqw2STMhWUMhUJjLlwvnL0r5XI48baeMHyzWnwUsi847wxzFj8SgJOM
1jFHuAAmDPUnjAUc0tFsPZt/BIL9GJ1kMC6VtJqhXUXd7qFmhEXLTF4vo+Ggp+cYdlK4on/G8kz8
/4C/8mBqwGY0a3ohYneyiyrvr1vUtaZWrdnENnIGcKL3N0mycwKzL/mVnp+oK2r2mSD95ES++Bnw
HmEAmg4/9hp5NaNqZWRZRf61SWnZkA9V9b3RfzUVuIt2VscO62fMeE4FBrzgmH+DsY7yBAtiNSWb
b9y6ihFi9mAyy9f3oJuySdvNOvCxz/jD28yGJox/OYImggeNzple3lWwySLGprfCuyqWkWqsevX6
zLIOoeD6v6hxPq7X6D647C6J3iAvz37Obp7fy1Dfwxy0dtFeRcK0Z6LP2V5s3uUPQIHd9W3c0U1T
IJJDbv9mLo7Z4hQEeY0iMlFOoG4v7E+WJ6omQ7pv+oUscyLmcdRFSrLkdA9vR06VGzbcJi+AV9md
sNivNH5S+X0ZPW0F6VqSkvl72g+fIit1iTo5UGSwnOuRM/OKkOK7KVm286HJxeTtxJEwQ3pZdil/
72BOqoHnC2xl2bJc1xf/97HdztZ2XPgzj2gDxL+Mri1LVFLnL4D9mp1orolGL8jEBUiNLyfmtsA3
a123+jZTN826AnKqV+wJSVnUWPhUhCpk0svx3+MwG03/AJVg32p5tuz/u/gLJOPuHvRzyi7qL9x0
w61k6Jj3sPrAxAhh2gcxf+QHxjoUUrn2z0MECAiT7mR+SQjCT/Xh++tqE8o2s+GPOJdWEb9dxsF7
J4/CGsFYScRktfp7rwqEGlK78HHcdHf2PaDILNMfPvlpd09Py1731D9KOANfG7IjF3Wo13Z9Kshb
qwNBz89busi8lgKSSpvW6pqW0WLVoVjAlawYLkjc0mcpJnTwqRRsO0Rs35ZesVcbH5peoG/kHnnX
KWaLO7W+ADznUM6TiAp+rOJKpMM8YZYxuBJnYr9nLtOSmN0C7bJ6trfybEtzy1m+97cp/azoOtkH
ScNphdXugfl9q8k5jK4R3DwCl02vQOn7mQUs2M5hLX1OCUmUIxKlIsx3TgL8l3/ktxZBwuYlqxti
7G7Jdjg2S6QMpxeYvpsAkyMDWpJtdw6N7/iqRzG/+vwMJXbLfs5U7Ipr1O7iW5WeL5vLB6hXLe2P
KxHzMwQhhDEa+oA/sewcFx2oF8kKgUqaY7yDc/DsSuJ/VqkRd5IVJVINOE/27SG/uqYU+dJPmVeS
nTFznt7JfEX1hLWTVIm7Hm8EQoBSe33YKuuDehhCAr4LP3x2c7C9nC1phrV67HPEpXxFEjRprrGu
nrQOBPFldJelW0Piqiy8MbJARk0a5cecigAkOzquaGvVGSAGvDXqGIWQPdNq3dZtRjG2UrP7TuI2
Fn+aaoR8vZCTwSKCpskc3VZdoLssYqg0WqcsElR762hAVPGrE7rucqzpFcE9Pw6JQ27KBYsoPzD5
BHEE3yFiG3Q9gXdEfynrJ2DwHwoyj1dLUq41v61ekN0GQ6DSBflYMcB1iB3WSYBG0h1A0A17pYpY
FqnRZTG/eObj064WFlITDw9ETZ9+X+iqJMljE87x5+NpyjzjRBtwjMOtJGXT+ytgfcn0KpCzqsKT
HvIsX0+INS34/oOSH9BN3Y3q+p3U+R8avmGaKAnojPoMY6yCxclzmTRpmWtCYJgeYAjUFPm2hpmi
TEaBtvqMOX+dId8/HQze5XbcYM3oguT5EA6EvAhQQtrnDhbu/LmUnCJRYPG63odOMs2w1nuJsxQg
AVdjIq+rNivBXFRm1nAqMv2q7xIn58+9VMJCEGMqMkJKm+Mh7564evMHoiSuawEEDxjeAQOCA0+E
J1DGa71LMFTaX02c8k1VlUcfA1P49WxRaU2mr1JZ08TQ338naDzv2ykJPmBojK8bSUjeM8gT6jsu
4p6RtWKsMzeYH+k5/wKHdfHhE4PF1Fyg9MiXE/q7Q89rp+7wq4ide957YaI/aNU7Ml9uQOQqfSHy
/oTNe2FqhB6O8bnRYCJ5BhLl1ivlCfMU+prFdCoD8RQaVNvVpSo3tzZ5ffQXCZsfBNif94Z5ttdy
8RSIwIhIva3WbyfsUaoXH3SNddbgnm0T+mRvKGDh63AUHOAwTh2kK/T/Beh5g613/mXqkOIRixxD
RzIixY7jagG47Uc7LJdgLE5nEx6MENdSdohsRJmWQQx62zlIN0Lxv59c2QBYFGFpggOXbstKNp/F
Pmn/02L27y9sgRwv4jo3bwds6yPeSoF1qUKCstODEFcEO+iipJOCawKZQ9no2cVVs5QDwM532gwU
KNDx5Q12/tf8N6hpMRNZeMleb5+GMTBWB5DpIIQ9RX/MfOKY/k4wE8LOZyiIL062kR01bF2lv5by
v9HMUV3sEGg6A/GUc9fKqRExx2ghn+54xtHoLqa+M5aOB1jmGL620WkhNYUUTyus7pUGevVqH1D4
lAp0qhQXPThNhckwHzciWm1NAjqK8Ke/VmNGg2td3PdriCAsn4JMqwdgfFBAJ/Aqqf5OQoJqzQN0
lvfHW5AMUHL6NmWg2zsin9QWbDOZjgNlgiF5if0UbGqtpimJfeJQ+bjhIdgetO7RYDOyy0oMiMbi
qnITz5HTJnFqJuNowUR6lB/Wppabdt1F3VWM/ajuTTU7FYBFagq1v8/ROOXTSzg2XDQIZDsY9YNz
z2Ud8xtG6CXQDdfcFWIFkBmW6i8WZVfnv7nJ3x89YVsSrvIcMrJtOxmlJIWl+rftRBYHNCLYnuof
sbxj02SQa7hY9UNnbtqHxhk5VQbxYaOqGZrV4xKhP1So2RK7oGMQyBPkN+KmKSn6PaHZ5tJUUvT7
eE+s6AT576Q6q7tqqO/p+6shckaWoJuG2I2wGfDwlPEJWOxR46AcgO6W2woV52meo2XKT+KWXKUH
OIwGAhKxiuH08hGC3A33EpkViLoN4Ih1qh1b9gVHRQHzVWouAlftH/n1EzbRS6ryE52zsgguvF3O
Nmqlhgu6SlMZrpAAlFQrSWbDgmHwHpmM1voLr2BaDeEDS1JHm4NRGxfGNz2YBR84BQkC4vj9NH4o
CbGslCcQqcgH1EGpNdGcdnaDxbaKbeeyqDuM/oDXZA6nxDLkKQ1ixtaJxDiImqXnaPIlPxomm6aS
yhYlYK3CJ8XUdlbGnydowEqPmUDou13U1FuCDeqmp7gb6iJ8yJd2G1gEj7rbwN5izOoJ1aflhNrV
0yEqc7qhbon5Y5nRrRu8X19uWl1i1sEovprhxprFQSCOTAW1/B9L+QP66g9VZ7qaBWVHmbz4qerO
t1K9NYIKEh2kc0AumYMh4si81N6dunP1yA06lXMW6d+txTrEYwHenV2ZKqze4VWlPRgqoCRa1QKC
3WkMWpDgB2/Axhse3MvBxQV7O+NdHpu2Ya1SFrsXKhszOEAKzUkfHkYvhtoaRblR+yiSDGKMlQ4P
bLzZNgiz7hoDITRF3lszLO3Ygw58z8FuSnUPKxO+yF94gDsc8PGDXW1bbskCQ+1YLkLrIBWTsR7Z
PlWj+DGqy4/62OGODjgkm2ztREW6kvMnK9nWbZjT++EDOz8hPcKfSMqqkJNf8q2U1EF0BmgCTuZX
HI9qwsLSVbkYulnP8orqZQtncp0haL0dOIJyeLB+UnTKFO8pK6NrKZGkdoNN27QP2ExegI15Swn8
jZV6YrL2dTVYCn6ahHKLpyQS9zpohFQobgATc4hKbTVtf9suLVmceDkuKDmR1bzEGYn6gd6PNuhL
YSdGZpfQ4qtYnoMjXXC7v04GfbmIHyKw15R34V3GOd7aL+HXV0qghZ67javrrucfJ444ViDigAL+
wRuSHkH941XvPb9yRlUd1J1yQKwzk/IkUYxEvn/ER72ASxn3jTJ7AKUAbQpoxWhK37qgASSUQ1jr
aLesEQRbgb57OPMnbfemvhGfgfzl+YpjPsN+n6jZVrBlyZmNudkN6dXJA8ma7WQvkW5NMtJopMMu
d/X47m8MFGCwrj8PaovFlmu5jb+a+OPwBtsw4p3A8PSwavUQBMypE0vQFI3kLoRfYbFY/XoC/WO0
FpiTLkErpgTFZ6zD9giBMCGFuCqUTMsz8vbxhlcxQ9VrZRLdzzGvRx+7tI6UEiy0QjBpJA8dSqom
O/QTNqT3dJPUODi9y1CaVUUCNZmhHQZzg0kNRf3U+mUVhi/9HHwYW/SsnplPbtEjmtAUccScwM3B
+BWzWpCLjFoCz/xqqgRzYTxvSfnfCNOo3L5gEj9f46sXq/16Uc9bAR5tCJ89VNNOC3RI0XeYC059
toSwcUA/uAImT9UN94bmiVMJfG2eQzJCLxsl+g6gdGvgPa6PW3KSUTgOZmLdrMx5jSScmcPD6w2F
ezzSEQYRyxaajanpDuZljIDHogxs9n+9c6WWeUSmCUGXG8N+rPlA3JvBr4bryIdzKA0b3jsmMMmC
16BDfaJTzBcSggdDo9JOOJCEmriNyfe4QjMO1ajGU7ajRXVxfqvAVaq3pnjtajqHS3JpamVNM5nk
V2LNH/f9wPkvrlBpd/PZqEF1d0oZTkbgYnfyZC1UUI/GoFgbiWTnlRX6aBx6Y4YTeqFng9ZDoXZm
TM3SRXalour1Ropp7fVhBEr2SGzPgg7VJNFnMrdEN1EAJD6lOb+B8WZIV/zh0U9bvVoZbWuqRgfo
rDv7zZIdUVNqcSF50YNJVUYWa9Ag1zsJT3zlkc1kHxtZrcwzjwrWUBubIH9nBPFWcP41LHFX61na
v7kGh5svo3ZF8VotzEOYzy2BXHVlfuqiMpYWSVcFG9w7c0rZ0d6yKHA96ES+D7m2I8EPBmIjBMVF
aPG2IXRYH1lkieaZaqDv4t0PMT9dEaWvp0uSjAgeAh4NkvLDa18XYWNjoZPef2clYXy597XE25uE
HJuHz5dB4V5cBuyOlAbtOK/3tHRKi500qUoyBBDvO1QTAc/cMbkJk9RvNhWLypszwdtqHmibVSB0
lxc3wHuPTY1V7zYHGjPcGX8mpAtwEonSey5mTgqLupGXtk1+eqpc1Wt7B7kJAYyJERCC8P513BIi
P/dnkLyJqwjamh8QLvKyvZumRAsLD5+4qByItZPQczi2UGo204833ekmVRt2U1H7EYIlsh2IdAL0
mgXSvOQ5+t/O2Wj0rNdOk8teaRwFhbOWmtw1UYkifiM8DG5VahWO5uMURy6gzEmEl7hx0TB1812Z
/Yd7DS6UCVCeQH6IH28fvL3IZrfjOFIyCVkZYsRTfM/FtJC6zMFi0zYTjPu0sHcfBj6UYS0lpmOW
ijbSCX/+HlDb93jewsxCLVA836fBCG4MrfLUmp673EaW55qLU+5R8y1OhVRhaJywFN2u3hZIUs13
x9N97BCVbNT6eayNiNF9JFWxIdqDUujRQBSOzhEmkXdbhJVL4K+D55gQ4dJi43Qv9mm6eEHpU+G4
UmXMyK9iiZhe5acqJpbKU0bM/Ak3qgs7zJdx0gGyOQnV2CZneRC53lqwoXxqLeQVUP2UEb0Y6lMB
VTUm/LYvvWFUY9PxxBZ+c88aWfTwOBb1UFQ0cITzgt3OdBvXS759KW2GTQhjWk8KMnINJKc1TO0D
B4OBk0keZtekiiIIMpPCmXUuYvjOXn3b38QCTKxG3Fh6gyfM+B+ZrJnOovXBVP6s01kLSnh6q5Ye
LE4mxBqkANPpBkA7f0PWDrb9ydVmtPro/DOYDkw0PtOSZJ0U6skbglkPcGA1wobczFcr+7O1/h53
keMmrFfkG9WXXejkmhgYeFLUn1AlPlTpHZVRHOzs91KxXLLSTkIzto0Tr7mrOeIhzbB6rdz1f/nR
dUwfgvJkrpQjgvFNv/v+vR0d9R6MlhcFx+XZoFaRNzr4RNUy8dzcaAVWgLKFn2sXaKgnDI46W4DV
Gn41KOmLg1XcGgPDyhPbyyo9dOgyRdJJm1Eo5l7P4+Ikr98rZoYIY/mqMBHzzKmJCYOTGLkDy+xy
YFKGltAmMiYZGfBHrKINWCOYt4V0+3wNYEJIDETic8sXqk+VeFO+nZPDotGBwQL1lltBk7zdXy7c
7jL7FQO/7lnztXW2wHxHsde10xLyQ9UnAkQDaUGycQQamCd7iKvC+ZTbzshBN5F9n/YVkQkfZIhs
5jmPPxq5jXWavVk5cnOXCUR5Ihb7VxGvsRMiyPacI7DIK67GffqP5deLzBA+z9+GxK4EbP1n36M5
ldnxjcwGRxT5FTgIyo8W16z+H+ZEo+6zGQAC7L0zp0opKWuPtxbNvTmKl6ymn6n1N9KOYi8sCmOL
zykUVgr6Fg+ANqyS7n9N267KHZhIfDCSxIz1nlQb8NIhE/XtX35+fKa1HggEpnzyI0Mj/qgvHOVP
xedN8iRiKXh2WCYCWmCJUpfIjbdDYEDrxW0HXF/RRCbTQSwRPj38J2MpOQTiu4pEbK+m/7P9Ezul
a780n5+881C6zCfSkMWHttFRhNRFQRIZSGrqVW0sixki2tH+X0vR/eGJRWxQxhyjACBru4K/RDEx
xVIJVpuxwo6TsI9thfDZqvYGUvo2vyN5XiZXtNWlfKUcrcwFh3jdICerjDt4SNvqGA7QFA9cFY3O
oprtVwRkLa1wSxY6bxYpWlcfIFaWrxNRsjyk+FQw5GchFBW1ynAZC9zn53y5Wij2nfx+qHWK+DOb
EpvXDKpJ6SmBuwHxoojxR9taSrNL+3vSW6Xxe9pEsraz8YdATmGopCDuRot+wehcC1Tc8rsxMpiu
JuAsaHWfQ+TziLQnnH6zY7gsse+CTnsojaqKwsQ1FisZQZhEx+3graSVpKZ5mVb0FgPQAAFyyCL2
OjLqeupK/qxW8xqTmPXgAq8vlmdlipqOnV6Ai/ijXuBaDe9nVKf4fAUbIYAtbmQdMIYBY0pn/lg6
7zzIFtI/Shs3mJ++U9xf8T7S1Y+ezTYNnHoX5P8X0s7n2uzJeSrtGbjANIEJZ6qAuwYjprOGFUmO
NcRxtjqATiseqC1Ip1KPF1bvW9U0MVeDfW/ozYaRqn8Tp6FGwTtseQKxezJxDUL/mmTudNvW/Mo6
USsYVLmgNwgsrJSY3fTcY7calUrfFmSgkVTkwbDrhJRso0k/N11pNo37AmQsFPEPNilLzuNuqu+Y
L/a3rPxm19Q6iOPUcBcIoEIIjZs+9vgws5LrJZNmRC3Mrr9tonMrObJCYcHIhLK8Opb+UGNzXOjw
wnn1Vu0FLu1hTlnx57QxLNZiJuf648BuNZuFZ2kQ2058a9XWFhTY/Y7NrKt7nD4EolSPoplmQeb0
C4KH12MFKUzTEja1q3R0etd8Bb16JX7W2WGD1sgMw9EI6ea3iTEHez5STi/H25y28e20KXNLgSZw
LCxR9bObteJ8E2D+6bvyZ3+q+JmCGr5Uo6tAgSMKdwfPXADuYUAQtdlPbtjm1EJ+Y11sO1CTDnNq
AnUenkFwIP8sFHmp7Ld0gHDmv2wUIKgXETSjLkUXnRG6A+ef4JOQn8cXZmMQp1rTJs9O5LekEuMP
U0CW0T05+oO7f5hEwFgAMepbGrUMgNK5Q38PUhoruTyT5ZoCtCqs/5Q/27y6Iq7g1Zal9pkQDwbL
qGjLx++7cz2hiF6PcVt9Ncoo5ywrsoYu+0t9HPd6GQyAv57yt96gkoETnm3arm3/J216UHcg1m6m
y/fJNQvM15PiDaIshhoOKNbcraqSwPA8bisJ1LFSDwwBfU2QhhwtgBMjIfSbMMHdnekWZ+uFaHxD
EfswY5XNDEiYdcetCezgoDBrgZs65RYDrwPQ6Ykl+jS4OSYBg63GffYnpWRM85Y71+IALXbSZNvC
GDz06JjTCKz6Ejt57vQHZXTT9f9wUNKEpSXPGA3y83hYQ3kMyH3qlOCvRYw5gL0n7fNJyNUPnoxS
5yUfefyxfhEMXoQWoWKTzyYDxtZphsc4qGGsW9sULnaKCaLpdQvHZO1Axar2B3ppsgxmrRdvtKrJ
bmkMR/Cxh/jtqG3PcIOy+5CISXIkEwlP7vXDJC3/NXWo15NqGX6NpptJyHd5BBN7rjRg1KBQNezA
KuSPt9qtNDS6yoppntuTRsyRZfOQUKNhG12J5tyVlWb4eSOFoiV8U4XgcsYTHTs0C0rALm08iS0u
OeRDI9TnzpPFKIi8A91w74GNvadhhsxUSjDVjaHKcLmcQlRjRbyIUgMZ0KhQ6Pq9OyqYIMtLgu1B
998SZrhVCfq0DBfPesFsklSVi9lMeqflIU5r5LZAUV3IhTjno4QHbxmcPTTgMGjOLd18Rj+ObteB
1iW3uXmiIEX03uEizrQOX2biJJeRtv/5biGlW1nh6B8zeMRTl6Bm9Ct9eGH49BTXn7EE+nrt7bUI
wmB2eB7AfztAgAYaslWyTFU8RTdDyBI10Od0TsOwvoJ6qjNzpcDXQ2E5ys4qkIPBiJojmtx3sK+H
sD96lAVFTs1x3wYWt2EBt9U++6jaS5vWCSsMi5go1SL0wmwLOm/mYl+m1lrzHjMimZlIRjqvbt64
tZikNUufzoYOOkf45ALKwUJFDxWJlAt2NxLDImeh/jGZYHLGkljHDHAnODL6Wo3ApXLDHKbPoEaq
xUP8+KYrZTndEdtv7Vixltjti0c4oiHp5yo6wfjGH1lA7BCRTlmadLOwSAk7Vq51U0fjLLFLVMsk
QDXQmejsB1+JrEPWW8LZUn8jnf0ly3SzvosdpE/5r0OVjdc1F8evMYNqvhVaIpkLcFU3Vk5MeyY0
XViYRgun+l8VnD7Zoipl4N+EumzwnaG6XSktPFsUXaGCrfM+9BDL5X9NLVU+vDBM9WDhMijELd9a
xgr9+qf2m7a6s2dDwvXhot97TCm9KjSrranNAGtWw8jjXtY3MovdppfdVDXnyR2sNTb4FKxBKJIl
Ru0EkCVQXYPSA8qciFmQXc3fGJuHrDWzLuT/GkudmVeVOvZDlLN1Ty3z62KzVOG/BmF8Jm2QFgW/
zFcw/5SS1RJbzqpviS5ECdxzWJ5fkBrRGlYzXHIfuzEiGm9MZBo21H9A8wbo/7+ParZRpk4quuaD
+IYomi+NVpiFFgFlQmrOffgqy2zcxSpyxnZaiesH5obbGlKmofWi2HLUAJMj1iYS1c/Jf21uaWq0
hk4e8ghSkQNfWyCu8SH1uOb6Zy360eX2Ht2m+5A5OzLqXnrKj4bEnQj9pjbyqI7w9nxXVO/q2YSJ
a9HBmRFrKADYxf8l5BkigHdUOsbyf22eVxZ9Yqq0V83sX7iXWpFYEjPqWkcM2J0NzoEbAUnFWbCE
CWa8/Ov/zUvWE63h8nwYpbQFoebiFOZ3uSx/wT1ob2XNE/y3x5CWXKus3/XOawHuoGxVKqayDV4h
cNjgEYuZJiQg5Gca7SxlvcOxeQkELgLSdilubIMIOK5mgN5I1oOJdxD49/kGDcUjpoUR+cRPC3Sq
pqruSZW8QB47ChBCYkVcd102Voz4lmdaTIQW9auQtVBwUSlzaAByayYZmBHXkoXNxO6hI0OYI+9v
bcsPxlYMCbc5sVyxwVewyivNX4az3rI50E98uRS6ulvCxoEY6/8jhoQmfLyrYShTMg4/5WeVONEg
RZyXxKfxLzP48LuQU/u1PzT3pzX6Um/FyaHzRTPXu4IkIQDF38IUrqmGv1DPse7MJ9FXNCJ2Wx/3
H/OliCq8KXhfRdO2h6uhq1pHlb1f491OyTbg/o0yQtwjdBaD+Fkfa6zOEU1LIhB6vNYVGmKpgqMx
LX0924H8hV+vwH50FQgEb2WB2f3S3AngqiO88ry1/0ddvlQmusRSr2Q4k+nEPgUJS7ISKmjfa5TO
jn4uPfKpfzmsBxpulEV1m0GPGNTAkBIfWCTiJTO4bsYQwQggCuOQ9PIPiFKQmuuW5YXgGBEmGhnZ
EY+3jokL/TLj3Mh2nOlwVN9885AroTHeBaGpIfOHb3Vo0q3xVwVhSYxOurehuB89GosF9Z0P7LuN
fsfPLCsJDLnrtmY+7ZvV+rTlUnWiW3pTNYIXdS2/mlKefFZeqmGVohPBHG7Hk7pcvZ8RHrFlBbwl
j9g6F1//WBwOcA4pev/QxY5/CLd1wazEhOIusZB0sC9Cox9SmqeWQP5WSfd5gk1KVIO4Ukzg0M1E
6kV8efgu8Q4CfuScLWqOx84F0BJPHMF1yKy41cOpQb6JgTe+Zxu/yMoJKKZyRelQq8nMUrz7UxA9
S/+hgRxzzTOjCkdwv8mBgrFPiKE9R2qS0zoEK2r963+ezFzFNRqrsJ9RXCZ8jTyw3Eo5LwQjgPeH
PeMnqFTcar69G3wMrTbKA6LAnbpoE/yEw//UQJgiquz+q86vZnakxFsPHu/CJp/F2gAW/EoJWAc8
QRkjsL6rHwSKkgFxImgLF9ksCQYXNGQQmVYCYeiZ6BuIO4O43NzF6rBcvqIrLV72EA9NG1vjeUfw
Xr3moFJzrxa7292x63eaq72LwtI4iEvtbGgUovVEF12iWhCJtKEr3OSJUrLOVfu8Y3IfREPXG0pG
j9MfaWU7zt8mnpWdvceJTWMJoP9bkzL75Z7HJMHFJrqQZMMMeWy56wAqinwSaqcJFT4n1lVQO8RQ
GIHJaNDB+54pdLTrS0HcrdLBJGulsAT69NH1sN82wLbKPL3umUXhbOLPezjGLIirqL7Oc9RT8pGt
YY7anGJrKnCBmxqUQQLFQutHzbfLYUL2m+3ls3Oa9AHUio/kpIQwft6R6SewDzYiM7iXM8Q7r2wV
rMYmjcyh3/JoMaESM7JSKv6u5Ptfl3D3pXsgPRIGjdRKz3x9PdKf4AA4G6hay//iduhGiyj5toZ3
yD4RsL65MAMoYCbhiiz8dYQT+cZwqc4Ryo8geMq2TEGs3aKP7b6Bzk1u6+3mki1nNm1fudxmovSk
927hSpqO3GmJbmGC9as9Ph1Zn+HMioTf8EOqqmz/2NYAciM+dlJ3cdxYKaXfGe7csXKZvE2xfeef
BkG8Bu/6qOn8rgUltJ8bFsh96d0lZVJ24NlU9kN0grOgDj1SPtOuswYuMpRtWE7PIBXJfFBXvytM
Ze4NecsLuUq1cyWj49rpDqJrksS3XM6Nw7KhIWQBu5PbDycMsOEK9urKXuh3qBd+inb+3t0p1XCC
SpD4HdvCV/9IxIeL4kyhdxxCVXLq8wc5zAFftT++VcPZC9pRWM6JmSSBiKn4DAoCHbHpGG+8VCzz
QBzGbW5NLVS6AHAqDwQ6mxPdAtNgIc5FNgbz7Y+Qb166uFfQSs+xfR//ggyJGnzgrS3sb+aekQHT
Qwyv9y3YbQt8/Z4EGX9PEQtAb7ZRLSYDByauUpRhAOyMfZsAKQyBPfTmpNTwkIny4FyvD/ZG1/AG
xJEG4t6FoKzl3fPEAni+f2JLHVo+j9EOFaj9WCT8b2lhsByHEGHFdVoX1b+YwZvG7tfFNEB71s8w
IGffgb/lANkEYY8W27/pnqkGaYeltzzjBmfg/FqovRZb6T6C0k3CULtcS+2UqlqdwLVlcDb/i3iq
imWnovZNQ4JS8v3ID46gMhrinfUjZ9HJ7Djd19fRl4Mibu1vvDZoXfIrRg53zezNXX6ZFqoLd9Sd
J4W5ekzYP6VFSZjMMpkYsfTB7RH3i6VnzdleMpIqAEmDrKfBL/gcWD0DV3VjnXHYSPQrFeI46PUM
viz8HxtmpWO0Y9B6bntK0lMOGoi6vhYRveKEmn3Y/lRQJEb0LgmdLruVs0W2xPVR7fcbNiOy+t6x
nWKzu8hjrtL7ItJIxGZIFlhj+nzBaj/rHom3JD7fR8CdSl3pImTHuhkGd7zfFHhNZozYmothQ8PX
g/o+VhjTHPrdwlbSW0VSElJUr5xnSaaaKBBrPq/5+CK71aJdIvL9z9hQJOEqLUKwAz3kneolTdJj
xNIJdpgf/ExGsRAcYnQZZQO65Kkmp0vxyBxq5C0BCE6Uf+Y8QKri2FDhwaslwiAV0ll5hnxH3zHc
385uwXi9QWE3rRMrD3aztBhySFoLeWYqVEDcizD9HDHi5r7LeEGHAM3KoIkosbmhMIZ8J6zBOkdO
kkciCcqnDCfct1LD6e17BoyN1juNTtEpOB/vBzd5bBYqUoEjs4SAmtcuCL+4qBPpRQrrCGb3b4Mp
UtOvZNnTZWk9vlBGLi0WBJc8/JejueOcGPev/k67+K3F9QkcAbzCR/W6kwz6QjmT65wy26t4ZNUO
QeQf2OM49JZghMmGEnv2hlGBUVBMxryVmb84zSO+HMWZXDpOcV2gln2+cjos9cwM2rM5MzHFc570
O6vTbQ9fJvHLW8QmFYLXohmwQZoz3MbL5jeYEY0hMit110kTIJm3O1NOLzdXbPUXfty+hr1uvtlU
0sifIWp1zFrKoA5+nd+YgbNkdiTdFKZoZmiQdIo6SjzDGDNE2Pzuk3Z4qNs5BS3c++dZk4PKPjy9
6I6S3Ev8fizDtdBAlHj5YdqctaLT+s3HLV9P3Fx/hqrmai4DDX++Dqu89ZZTsx9xJrfysmW10QQW
rRgN5NFffE7wmOVldKDkYYOboE5UXOT4xYgZbeKXD/lTr7tvcl4n0F8axW2CqROlQ4rBQhc8llXL
z+JDNGx3CXx9hUMDd11Uwpd10qV7zbayi+7Gj6aMAPLQJC1Z5xPXMc3kezb/nT3GK7rEzVFbRXjp
Z6VH76jc91pk3e6MHvTCrpOUTIZ+QlcAhcWZcee5z3FPXXLPtpz4in5W/bw7+VqmGKdvhl/EnE5S
RcuuX0s1o3iYAsiIkTR0zOV35z5ZHmKeifLwA1CnDPGvjaSpn0rn9AcTO8rGnkzRa9twZzBqnXSJ
2sLxnfHbiWAylzm9Gz2facjtcY/aPdLnbJZ9jv1Csue+YF1dLKGXO3FHc32bC+PLUzAOhojjRr4Z
cRP6OW1sRZKCXJ++s1p7E/FHYGOQ46eIiM4QfreS1Ne7IE/1N1v9Th2CjkAAGwKtttLm929ohkfG
GLc/NdYeVt813ExkmXKyZgAystVuW79Hp5p76vFA6xRTX5luQOWQUlN2giIgYfrqb9WHITPqhQL+
ZlP2zaP3pKy1Fo95Uuxj9pQVKMjHPAR0VClQY8Ho7EOHdns5CGYG85cnCBmsCGIaL52QjH4Zusng
jiqlxtLCJyvcGu11N1+AaEi5yhpWJ+W7jmyH+b8U5nEmYBOQwLkSlYSwZeYB7Sk7WS7rvrUtzaue
Y4N61Ds3UbvoqnQw3EVjlr+1wZkGvXbQ/rZFnU1ZJJ6PGfDDUN6ApUV/JCF+PwwjVxbyoNB47eWl
dbwC/dNzNnPN+/Ld7OMNzrnmavCbbkhad0pmeg3JsRzkomrjoHnWLBAkJNm1VMWn2SU3Eo95RpeW
Q1dltcsq45HdT2i/yvf4CRw4HI3AHbEpaki+wf6Df10JQSWXX8oYNtv1QXAC8i/QcLTJjH9e21V4
XF6MTnGtF2keguwYa3d8URI/4BU2LuK293xxtliMQ4pqG2j7HdhhziZPut8Sz/wimJROaP4gRWY1
egWXrWush2biHI9JXKtBVueHcy2obWB8S3LT7o4tSI2W8VfOBDjNdm2GlIl0XYBsKw/Uvho2eWhp
F9/HAAzrxABok/94dYp9AwJHj/hA1GVVcvFAOptiIAUdyfdn8R7Ha7jSXdB9coERA3hsAt8CXhia
ZghwOPT1oNqJ2rXFbP2zUUJwlAf6YydPCyF9ackPb0+c1OEQI9rcb7QDMqu1Ivw0XqJlo4fAhpBG
vZvNTHWArBnLBVWGYYs2C19y+5dYEv/tQDeMsUli6GxkSrKzz5U7yqBpilOCI0IjdteGFWODY3tM
4AHCrnvCBssiELKSB1kKz/JbMbxPuVh96X0cyKHgmDm9Fbl9pafwPQMQhrWoi0SPqHqdBO2VGJGl
CfqtKuD7v+AUP1D2ESEkESegVEHKvsxrKSCrPIbwdDI11R+m4z16KfJdGyR3aJNaV7DL1QXgXyLD
9qji7KfPTz0pJuEHM2XQCub4K1qGvU5biTVpFBMMKm+uI4lqd9c7hHF2g4fsJCAuCTV4josYCMRv
xeEFgxEhSqQ9xMAaYsv0lMjKBcExlHjzgxhya4egzGd8fsnH06qcoDjl5YhsU6cuMM9jEuvCmKCe
7t31rmy851YaW281xdhRHVmJJ4qWLEar0PQ1z/qv0/fmkVp1lRib93+/nlqg28qYov5LuELOdjCf
E2JsP21aDxM3mBQT6HOiUa93YXbXQ25as+iI6YeWo32Q9YNmp6SOYDsUy1KdjeLIfSA1JAubGAcs
M4gyENwrsE4NaCR+13JonAkAjgDMy1M+2w1Ps6X6LkRgbPls0CaVe7wBa92zJI8iSDo5e0PCPTuG
S0OS4Zzp60gWnCzvEqGV7jmNG5751Ol1GU5pKiDog07mw2o4yLwt4EboHYYrGYmHBAqYxsSOjnJg
GU0piLvGDXLO+q6ZZf/lTuZ2kMhDlAOVhIwuZniS4kJJTnNZgJXROTSrIioMr0Xn3HELKZ2LOGNj
8hs2kuUY/F26llU+73xx8ehfVsHStsv3TdqZMu0QPqJTCenZ9yINyq+FN5OK6rj++Nm8Sn2nvxKU
6hmEIli6kpWiSqD7wfh3S72/rFRqUowm8/ED3OBnbrRFbWXi1Ut0Vk6/69oxO6KhWmeRTcC3FnPj
M5wHTIakf3SLV54SQ4mnsG8qCL4qCMRVH3RiDlejC+2JqWir+WFrz5MxAjSkRo+uopPY4z8KIIOC
3yTQIEzC0BvHLFbib3xHHm9NSp+WavVmWOHpaXNHAE8S6U5n3/1XjtnEWm9+z1Mmd9Bp7pROVYTV
SyG3Gae9G9NKhawBkh9grimkvBK4xDNwEwE8Q9Kd2EQSMkdZ7WibzDUsn3i2rqJeJi3uJchPC/4b
ESHISMArsG0DqvlRtoCpA+GAtpbjf2IdlYuprkazI2E8+ZWwiIpzg/OzlkPYWFKqoWsOB74akzJD
8moqDH/c2gXqOd+R37zGH/hwd8XFsVI/GrXGGqCvVa+iXRRtFaWY5TqdQesrLzbHnWkUl6hJJcZV
DW6jiyTPII+7H1nhrx5xj7nd3ql+8fk3YhQikmTC3UTNMOhzPDYx+CFKZHzRXhObB7Yj7VcmS0nm
2/fyStCSIosd6dJ8YRNIl2vZlRwb+OQMHBJbmIy8WI5dmhl7p/h2JJwaVR9fCX/Ixe2xMJdKfMnc
2IiJbVKrPoIRQVVASYXfK/W4V/GVebi0gcH6eXV7LNRpZRv86SHl+3AqkcoXJWhiWyG4q5Pm2XXI
gsVpBTXheALELNKLNITD35CfsJN1HBzybRdceP0z1XvihjYWFhjUDTQa3fMTim9wgyuZA9y1Pphs
YzX6LQpfztLtz8fiAKQFbzRbwjSsTsX41OGMfzJcYZrkFCTqFzn38ND2RNSGjOluxj8BG/tB1dFu
jVWUYqLRM6EsS6l0TOnoqHu6SphwkBCFiNIMQiTgT30eBcoID+LX7Xc+8iiQIOzYuv4QDf7rJN7X
7lezyADEtqHRozI5enO4q+qzu+g/ieMMt9xNX4kasWZ34TGJ0iWd1nc7jDYC6zELlDg7R6KGPX3A
1JnIgdJMMcdCGmv/f3vr/tamvMt/r3rbtqX4hAY5ZxvVxpvgQxF0k0SoWBfH1+4TsrhPwseJLNL3
vmpAVs6SwFy/Wkq2DYFzeTpGQzukJHvEpvj8NaHeuWSBkT+1GWl/4rSCbUxRVoXzEC170KlrIVAC
irXBzvkVVk4cx1Nd9SRxd75dgD57IhK+uVB1LtaCr3FdwFLpP6wW7hq07bLrCR2N61LgPZX4Gjhu
EaG/OD1BCJp8pAMGeXVsppeI8yv5W0qd98jT1Fl1iphEAH31Bt2JpENqjn8L88O2uq7oXPT1flXe
6WG34zgpYl+kCImc0VRuPUl3v8I6fItlgtIQShqRLhaEQEPF2quGE2UyOYg6cWk9veyA+1PPaSAS
62D5V39zq7DDB4quTXi2N9YooX1RgUs3I6CdPBANkg23KrtrHnslH9JSqfm7z6cqtIQupI6mhKr9
9+zKoi0WxUHJrCVgLO+QZuvKcfqm+cYJgQWAGBb5ogetp10b5hTrmpGX9Fq7n3tfUqll+PuTepd+
bd/aU6Z/MWRJa/PLgQfIabpyvQdKRDRnLH7TNi5dpkmWHTX9G83FGBx/P7GXwSj+Nmsj2YzzlYmA
NZwpv4cdqRF2hbO6WUt223XuIwPWo9BjKy5KJy04WRyoN7bzeQIkuHCVNQ5IqVYusuYScdkRUY7I
zsz64B92KBW26tS3y0q5OJoAxvvSXJnheDUrqjnqNPNOI2cIvtBJGCQk/8HJe/S6D0MayzH2Kjk9
iQ0hQUhBEYs/FlXzo+fk6WVdDKDIUdNiH1fs2kVhfhZ56CpnMbP4EKL7IPQNxYQxZti0VBM8vH7z
zfRKAGvdB8WxkiZE1XgGvnOtJwFk99DypZ7iWyZPzzkghP/S+6BP4iZ0Jhsum+EVBdvTyp1wzTm1
VKJBIcBD1ZDgAjDTMQO9M7ccw4bbU0Bs4C1fgpkkY6lJYWMFaHaXKuEz+jcHZCAFCFKUhzFIozJg
OewJe+Y6XA6uNEDGdrITb3wuf+S8lMDTnB+/WWzgZYwNPAzHnHldA+1LAxotXqnJscE5unTysFD1
u9oe4r+del2p5caZUvEdhAYAtUKTUIF06G1o76bKFra7Rly03VnH8sW+fBNn/8cXZ5WrHJ7a744K
un3Hoc7zWKwWIOmFKDEdxeblzu9WN1x2ps0w2oRFYRrUrdT+KNjqH2ZWfn6POdADjSyKPHr29SjR
J+zcgvxvWAyCDtql9h8n5XFktHqJeqC5nQkyKR0h1eNsKZYXZHR3isYVVXK18nWMMi4qK74qwy0C
hO15vUDeDgyWBqIy0JfAPr7SKfxq42I2npQSTbvuqqFEOn84IzrilH5+sqrJim+vOzWVCv+sTAhc
7QFfyC7QNlDV0CpbO32vnAUuWPlCERkzXpDcs/2fMGJCZbZ/zh51dUnyIcILniq8bskpZYfzuaTj
mtzcxStzDdCPRPDsNi2WoJUr3hnevmvLI+XD6kY1nWJv3W5zhrHPUL0X658Xra1XTlzd6bof91O3
vEvTXe2RY6iMEbDAd0TolbwhHWtFRabe8lXLbTPrUzh4KZJCLpgI1e/XfOCdGG8R1LjZ33k9ILsd
6gnQk6XwzHzdAY6pF1ygRqLwSz3ff0lxuaFLlT3rmUsUwHJFEyCwZX612WmWm48Y3OPNKrYmJPAH
TNrJWKWByAV9dV5DWQ4daWdW6tgRPK6kJIoZzGhFWPVGO9BSRoG9jWcxHycSYiQBZwC4qU0qGZuL
JAv9Ux+20xebYuR5DjN9+UpCFl8+ILVfYE5zQunLC2c3ZK0MWGmP32o0MbEWmEz9XM7xognvvanh
Q3bXDOdvyZFbTw0eb+Cb8SDmxbP2DmIxPyjnBZLqGYki2I1GBQQD4B7brE0wjWZgkL2Huq4QIHBo
pRGXMRgGJP2ZAJOrxWm/VfMqUORS8rC4LHuFqBSS4Ps0gMJa9KFMFZ9I7dArEbOJVXZE+t+ICLZp
a/N7M9j11d7H24TfzNRpJwobzzrhliyaGMmiT825KJuVGxWS/699SfQui67FZUaIpXWBPPkk83vX
WkP90D1Q9oTelQfgQOEjD162RgNoPKKSpNXzrAAEQTf/TgbK21dPztweuPJsLVhPKtoYcL3/O4uw
w8sYFcOSd+u5462t2mp6LN9nVSGYm7m2LFHIOmqkKoklCcnjqauQNblQYDx8JzI7Joe5NOjvmWEs
Nub79XgVHxYo4S0O7UVkE1m+3pJf4qltZUfO0nX5dvLKxMKiquEQ5LONraZwqzRfVLo/q4tHWeSU
Vt4S8oZwjW361w0uPbqCEkA0d0hbP+eECJ7SUC6JnonErKSwQ2ivZQCvefugnrAwTC8fo1gpz7JO
NE/kbsxsKciH9xUxLqd9NlfAOxipEIWrNKgfVUnL9po3mZqIpDBOSFurma+dQvNL1Evv6Epgt1wA
x6m54MqwLjG2uHX1fW1XEWIY0jCg1/WQUlijR86+gRtKzE+DFFtpHHzBTGL6FT2aLfyq8yMLW3cd
f2nTK77Xu1paygdZlHaD1ldjWMJQnk73FmIVoKmB3A4r68xAI3BNI+qt8vTWvDet1QF8m7Z+EWOi
ZzDPQ9nN1yAbcXWiBvGhlDsF5mefZJqwN1ZubZwIb+GVLqJixwi4Lb8mjTBIRydP7dXXAUZRcaN6
8orfJalUDji+Tvqk1OsbP5Btk72Nnk8HzD6kQEU0rFGkXeoa8A38wQ0JizpX89L4Csq+YrM+3vLi
gNAVIKfbUqSXQDxtC4+9BjXEiV3ODG6SrHzSVY05kdAlToLt8Lp00AWGfR+GwAGUGK2JayzCIIoi
zQVOzRUpd0qKQsiQEn9BpIBB97LJ6XIyCuW1MHkSdQKYKmqSq1wCQ6AfEP3WRtjo8YVTgjglBOuQ
m1B87a312nLmay+K7sjP84+GMbrQtKePpcpl/u+jr4nYklEQqq4RfNd3k5MS+LgPWpjqjEac6VGs
hOeLxDHU37U+4ZqLHmKdwno9o0hu6tFpXHE5u0LMk6j9Evn6LvBc6mv176XGPvqqU85C5DDubKgB
PvM97eMG5q2QLJxciRD8L8fp33viMF5kKBoPVHK/nBI6yATp1BUP/RcXH9ZM5H3TXdYDXcP7Msbl
AV+J3G5WGynJ0AcGq07gJ6ca8YJITS6vB/Z5v5cmEuio+k+2g7e1bRmn/RHc8oxzM/2aYUo2WIBj
dMwE2HVjCoL+APVjTcraHL/zlCSVXDxNwIjLeXjFfZ/RzqaZNFwe46r/PLl0htpQTlVWqjTrVbm0
N3qmDNfx6klsfoHyUhy7rbbB8yRRxDS64M2XK86F/8C3/O10DZDHZ22FlXmwtEXBRQN445NspI5b
Cx+rQPy09WxbNtXvy6+t32PliOdgEexro72CENp1uFCu+lLy60Adv8NQpe0+9rmqM864rbdCPs6M
6fIozDo7g0Rrj8xc7P7CVDFpj58E7Wx4YCOyEUAmqSBKphO2P1o/hrVHJIXj43SkQmBx8oNLluJB
QVbS7g1zITDmJUVUqRSSWbGDAz2oYBOgJYcGsH88tM6GDnj4IZ5IoKDQMVGYNqvAaTqhbO9BLwln
TvSNu3wJC2bixnQFLj4/K1kVpVJlwv2J7zsMwcgqhckYvgx7PR5JWR2AIF07AhWIG6REhsuiuBiA
PYCivtvtzEd/1fdq87lvOk4PbczYKfghM3X02Y0tyyimaP59Obl+UD0ZPU9COtyxXmkJZ0ZumKbp
UXI4JvLyhMuxmAjFEJcr1mEIisP3fPGMllUiB+J4RjEKzQfwSXNc9kjNe3Xidy5TtQ4DSM7lfuOT
eRmTul66ddN+2DHiMYbCDZgkb8Afevgb+5LNYm8B3ZDe2a39F3WPphL65dgNq4K0H1j2hW+5GqkH
YDS3mM0UHXReRsO9cCxOfDaHudWYCJF4viXp7P8D/FrHzAveseuAPEpOaGNXWcF19uFrTm+D7Pkd
90x3U7qldFPh/6hHtppk3t+2nDMCzycQfkzrGqz1d0Z2/o2GKpC8RZayUWB/73vGOgWYKmyZjN8p
f3gK3UhkW81dxzmXtesULNl8p0zvmocZvK2gh4pTxfvPLvkRUb8yF6xT6SYmaawvZbEqEdme8WSt
qgfK54ZIPsmorhCKp5GxgX+zgeCSVsusm/JP9qTitB9opan00LQbLmJU8o77O01W7t1+EoIgJMJY
tf/3dn/O1xHm20/sHb063XEo7KfMnYtgcmBL6ueGHK4gBh73/aFwxHKOdTH4LgOVC3QH9QlhTsE0
rr8/+wQMID20V9qPo5goxMb4O70PF4XmP8dlL11EbWQXb8MAjBKxwZhqtPuGI6x4KMdzYrGUzpPB
HgF0iZJrg4MFIDPR7diOezuxAspxF0xuDsZSh85nbmAbouHFQ5lLiHwsJ7DW9A5ad9bjvo0Xlqnk
14RltY8S1eVKSZT0tpTTO6Ciausd468Ng+IRfX32uI07/+exJaBcA1fkJyeBLOZPfAQeTAVaYBnJ
QDcOu/oyZQVSexGSrOMBNUTWXeYLOo7symSAaTEduHVxereDKPQ5yC8lIqNe/eT45NoM1SJ6ZkNs
W9m0F0oe4tSA/lzahZqcOHZqIIgAiCkZIBeZER/+5LyrtaM9UO9mSaguFJ3oToUW+mz+5p6hz3Dd
bQyz62B2ffezqvkVAwMOJHTl/RYszF9XLlWbedJgelJsoFe/TpgoEYJAmPhSyirvG++51zf89RNn
JcGwnmJGh6ipBnrgPZmCsp5mEALMfFr5GYkjcoKm0uqAr3ulbucpjuUmarbj4JVO8sOF2I95SiKu
xmz48qpLN+qBKXp9GovBUsiCi2RKITGFcLrq71E73pDcyAYJKzEGP7W0aa+NkQ4uK0AZK1eeExbb
HfqZZHO+RqYNoK1jv/n0NtQT8CSbc9uOxFYVXzMEGBYHfN9O2pd5k5M+H1CFAFChxW8fQKSAGnhS
iNEBcIZJ2eYGRk86VJBhPebmaLWY3gFtV3Pvb2Sj9N3O2ulZ8iGa0+cNOsWHGYJCAgTq/D3PjJak
FfY+al15S+Jhqa0An30oz5udNxEJjZI0bSy8VcwDjT3WoLULf0mgyWzzvkF0VzlFjrbXfrO8a3uu
1sgaCtv19d2JFTCN37RI4Vw1A/l6/jQ+JhEiUXSm6NuTX9WvlWvqMzo9bev1wRsOiR6JCDND/e2c
u1icCuQlqHPGaydLR4Ch0mLYCgAThp7qkJDAN/FUsrL2ZSw1gMVhLPRkuFdmWwFYeL+xjj5jldH8
WUDcMTLmFTeU1l8t/XuzpzQ+eatX8d1RuEPEnumRen68m5hX1GYCjC2eKd1nQyQ3d/QTYJX/b0Cj
hlx5nprWpQzeHA3lRLOQgAYVWNhOx4UVtg2YiRO3/T9dfXTGbHNzxlvz8aAff+eJei2W+IhzpH59
qJhsxHyuHiM5jOrKNZ15Umv/dx7LMsJhjlvRN+lPkUJBrZ0X6HF57vo8hMCfJ6G6BRzo3R8FKca0
9FPm+d+2r6OARvjtUWhKiGbYOXLQGwXbX418GVBjg/NXjO6nOCIgLDjPVLsoVTze67OkmUUchEo9
W/Kb6gmUABsjxOIwKiPxhnc9ezB1LBJf4GA3xPAHQHz0aBfxLTqdeN87WOTV1i1iDab+ju+9+U3Q
ozcrXiYN9Ou3GEWlgzMl3hPH8HcAfkw9e+7EWJXV07J0UzhyPOG34eNW97Uco1VoLyUUo6zcphak
BiV7jTIUi+M7WIiQ/X5RAHBHnTyUpluZkSAvcBVENeiLxtnJdi6sDPjPsem6jN9Ii5wg7tJll/os
UcmbGiiH71decWQWDB9GlzRYQPyuX+EYj0+YHHileZcYpHGeZXXzkvYhUWqcP9MWS7JYELV4GBEM
YMaIwsm7NvC5NWw3p3i9vvrl2M7UWnYW9tf75dFlQtgHc76/SrGz58iS5tXj3FnU7XnT0fOudxFT
29Ek60OutOWfvnfpmXqZRENKRt+aWN0IU5Pbdua5MQVkDQSTDGHBy7+GJ8R7Nhr2UE65HKlDsA5w
/BsrNKTkTDNyYSmWZxQRMIASL2p/6Km0TqqeH3cNqtTRSGZtJNqQrtnVa79/OvFO1enDCtM92fW0
j6EqqLMpT1Z1jCQhKuFLFvIfvOo12RCacMEbnNw/qqSh+wCEdNuFjVEEEBnq/Mhwre2uPTQhc9TW
jeVDOgHSEckBi/K868kRplP+K4kYKeGOs6huQlAgnU2I3dcdskFRg0XPALnOCUV+IcDCI6RVTTI1
XRjoLWHVEkd5JZbibXd+Z6EiHrJjDOutmnF32RlRjP2gFyBTMZi6Q7iod2GhOE7xFohYxnJO+eRv
H9dvuZ9MTJ33VcNG0dK+Bj7S/26g/EowuojDmfQcxK6byyyXm+VTn5an/LrPeKae04QROOJ+vCEa
vrDREGK8WbNcbn8jY7IT/Fxikay47LN+AWj08J5hPQSMyK8D3ptzCp9w9F7twcbDq4foWVJPei5F
oL31ONLFBmy7Kvu3tFJdA7quwnd3NC2zhe3IePogzYxJHlOO6e0eeXcVnbtwZwGUpbkRp0iHkLKW
LqOVHnoeXKGiEExESrzi2wSFLfApLE42X8frdf8GmcaB3/BOZJ+XP/fzUbZDMd8WJyUFjEfKrdlr
G+u436m/4J61oT847zkJbRz//yIzH1dqCG5Skj2GtSSgBuAOm+XSsGRj0shfC5bQ4lWj3/sj9rKt
+PL3N4cekgIsoj1Vaf7TurvERJfwwFKzjtab4mspf30EZqS98yeLStFaoDW6HlRiYlobkazJYDbL
BI1SS5bAgSAT+WhX81bXdJ/hYcvo1JxZfXxX/kH5qGIjCmAkXUTDQ2Tt8eGJkd0ORuAB+hS3/C5x
qMRZ92JXPMgqpOWkaQuLuaAtMnUJWbvtIKnzSkUTEjH6I9uzsu3Yq7Iv5pSAQkFG6jm1IVo+x+Jj
N4N4psM6dIav0ehSi0q8+vzGnTP78yiSBBUgqCfPDqqfzFTjbrEw9El+CO+LqhOhiwmoNFTNO9Rb
uARmAHqXuMFR096xdjWm1/sR/4wmnPmqAhK58N4Lciiq9K93iIyG1JcEjWAFOwwxhRbpxR6VyrKy
mdvzJq1igG4hfGXfqig2qiDLicIKyW/uDVdYKjY/Oqk3BxGLcqSMZPoPkIERT70q+5ENUDavLWsI
ihPWThLgXzOUvwM4G81ayK7IzXGQ074C4ndNJ43753DAL7xzwHylYSHb1tywjbG1W2FucNgqwGyX
4fk2PPH1Awcwxb9E4yPr8Mf4G94+dn31Lx83Xz7PQOW/wyEJuWvnCDsC8+I0Ds9yveXe7t5DydIU
6IPL4LXwShktAnp79+lS8OvVv3omindecELjX0qxNIOSVbtj4Ry9+0f5jdvK+fxwC3kvYqPbQ52e
v5PcNag+reMPM9fLF3YbTykuxEQhF3RWncP9Y3qpyDB/m+0jLzG4Iy8NCyVbwOLey5rf+XXxGdAz
u02kSRwPQ8W/wWI+t9jd1LxGgEtWyYru2LNq1HHCTw9TK8FXdVQNfSgS+GnEZMheFZ5lN7Z7Q4Z5
NnlBQfyaqi9I7JA0pOcNuLwG4Y1Gn+X/5O++6wz29eNxEIvvc5NVYrRCQpIPZ8e6pUzjpJcwhnYy
P4wkSyQeX/tKCIpMYY/YaWx6vterT6VWv1MIeVphArla8zDVp1AU7rLtYJNwe37niFT5ZeSUGPYD
F57qJBBxJF18MN7Mz+FXCKpW/hid6AryaV7v7Ec59dwuJoDQ7kbZtzMIWztPqZ9sxqbftEevZpcI
zcTM8eMlB9N1h/GheccQFInN+vBS4Nnc9xXWW+UAzjmzATAI/LQaNeNYuJeemt0c+ZlMEErMtqmR
fIZxVElsapG2bwlUfqcb3bthi/rko/66rWApuSYV8CAGE+yixYLE4fG7vQtB2pXFF5NSvx0pzRJN
Kg0jSTi19ZPXWWDvlWEEMydlDTZB1L97bo4hmqWCldvX2uMmWXUqaBAhrDFkDf5DCWJvGfLc+PiI
fJU+GR5k2twfklMGoDe2neZJqW84Q2HVWtzdi8RVLhCwOs6e6n/ns/IKYN2sX4oTyXn7RalcnIhy
bP6t/69hXOzTtEV4yrSaP3TLS+kikj+hDpuZY3xLMU8R6W8WFqpMAg8A7AHoFFbRLEPN2YAwB6pR
Ets52JZQduLBLl0Uqd4+r3n+2kJAT6vT8Mo9W83s5TkxZ+fxsyfYSZeYMckvYi3alkisDHYrw8kT
XsDfCY46DHHS6ohQGbheR9NPXzBO5ETRj68vH9SUzKknkNDGAw1z2+DzfxMdivkIHr4gO/uSSnca
qzWHuOpRGeaMHozyRbUF5Q5xdzR68JR4gElwEthbmg0pwfDdT2/eNW2rmlyXMRAxFNgJUbJkP0lC
vp6qXt0GCvSIF2Aae1OX8Uk1RPTvou9C678VbD9KL8d780ZmjeUOXcF5kbJhfdSrFvYswgdWqno+
QnLE27hDaYqsRTW5lx1+Fc2iNIbZUeqa0d5C60QekmLjSNYInxa/1J5FHiELDZNc2q6hhprV91rN
f+WiFQcATaIoU5xF8+SDXJwpang8oz1ECk/6Zd5MXv1AJUX4DqnoVeQ9tZ32LAMj0Rug8nwCQPzk
L4MoPSacKlDHEbVYOqxW1/ASeqJNOrr9/VL+9K/Bo7ncZOPr/1meRzm4k3d3sQ1rS8pjGwhdcNRE
rG3TUqfNISva0USJXaxGrkavWNGXptLpvjj2RSkrG+HWrUPkjhkS9wT/gAJ/xLjTkcw9FmyZanrx
m3wW0gygzuKkzRHf23aqXq5sriOxhsSoBioWyELbfA2FgLnFLqMKpCYnC87NcpImY//InSkYPmsz
cVmfj+CBWXy9roUogK727PRoSWNomfenjI8PsBjZ2oRIoAYlaXxtaJ5cUQz/G20/IGn52IsE5VJp
iD/oXMdNCiPKjkI/qJB1CPGnFsVNHipBPrsS7gS4/k4Gqw13rVgITnxDO00HrBFM96auwb3ivd5z
4Y2JT2xk+qDHTaKiNQXJ9GOK37k9ZAG29xm3LNwYeeYD/VW/UBAUYZFBiuEfyx5CrVfL+ie5BTvm
c93lVXuV7Bd1DCK/Gd4R3odBdCfTXcBz7h/sTmumRAmqjsADNj/0DGPOtVBc2EHs1xCg9xozMA9A
Jmzn+L96kMZA97FCa1k3Ek9Y3ynGTeJjzA7rt7Q7oMoP59MAu8NNiVqL9DfkWArJh4r0joAqBB8E
K8P/9BVCRnnx7qWG160k0IFyve+8KAuvBroailGDcz+M9gF6hIuwS4wr+8mlgYC/ewn9TVWdEEde
Rthmg1EArOqMDfCkHEG3LN4YeuBc99mqcNSiAH2tMkta0Mr+Wpa+RYoBRX4c5V4tX3KwEl3IZBMr
SPbOWFg3JptT5Tawg7WXbsLtwOsxdM69RuEhSdWRb79VjwZH9njiYrLW5pPU46ZIEPWzrF8QnjnG
TdjyPWfUu5QsfIkfXWX8hI9YeFx/vIIX9nI43mGacCzqy8KA7VkRdqoLUmAUlHop5Xw8OxGWwuQb
HQORWVilxN4ZlUmlqkoo0ZZnuMR3cSpAJ2+N688SOSyXyUqpwsGtRKpe4UaMFMBB9Mdf8lLkJ8NM
ISfU8jnvWd/VSoRBzAN9nx8YeejKoVSQu+VnYTy0doQ1jx/5vLhVr9Ou8oJ06QtAuYVWjwIru2Da
2uHdV105+5P9Br7ZlZXhSH30Xgl2pPYlILqN1r1PpWu13AmI2JzTCGrgUKyL/WycQ+RcGLmN5Uiw
Ojf04lH0d7hZU7zuM9AvLG6mM3m3VPKrrnQ/5HP2/J30Mg+CiS9TRQbkl1y2Z4e66XFDI8SfGKfY
ZKmFL4QdQS2wUQYftR2Dsrb0Jgb7RTudkX/4GAhCCvo4Ia6yzdgynorNqibLe3paW4hIYMD5GZRT
94mC5/sxJV2eKufgTwaX3SWqrqyNhsfvUlaOv1fRgqIPZ9UrijbIVwZA7o/veb1jOMXWAAI4jv95
Met9DwITmUmOxO43c8w2wwdbKK51TeZMvYAwhZCL5U0+vAfu801HCO0f66cO2AzO/rGXzFC7Hhkh
dx7n3b4BLbdvlsjlXxxuubs8s+ryjawf9AF9KrCc0tVl+WUFw68ijTDNMeBBySsOUtxcG4ECl4EC
2Xbbl1GZrqOJrxc8DV50BPJpUq5HYpReRJsbMb6eWF1pZ1j6p1HSSDK4jzepnDumLhJJkeBZfqGN
3p4Y8WJQQYeYgjDhIhQNy1hMyztq8erD3drhpfxI5oETFTz8QAA4bX/1jIrRbIDoHGYI5/8ITIHQ
6xEw829L4V+MTa+KZHs2hmxU3nMs/dlM2zXp06fWc42jIdHRXB6JS8kGW7sdAO8zmYMtrzIRLI0b
eiLXlSZ2nwCojSl+3Ur0Wc5V7pWjUza0aAn+JHlcxVv5QoiNNq+wpyPvqt71hmMITM51tymfgLfo
KxAKkGvg7kV5xz4VMxXN/pgHlN2C+7EOisi0wzQ/J8t43RCyazOZrZFXCh1hhFr8BrvgxXyWiaye
DwCVbz7AguZvZLQthyx+YKfdoTJzzXTszpXc+erKSleYmnCnZt4R9IEbFFq2ymMnjUKxtqqXpS2X
NdWNlKfqHCHjlS8Xi2K13kpua7mn/29reyTtSnuvXHpfCO6dXVbfYyqOkS9dryvXiFfyVUMKATub
TK/ItNWX3Qgdlx6MZD5C0lB5pwQYqWcfY53t+PlnBzHWl2ODNIQxPjRrpAu9vJPyKq2CENBsxBLw
TwY7xh5EYzVfC9qd3VFTopF5xie1bRyCnsL3qLTlOV/Lc/f2sdEIYrGOzAsDkI67VRAnnzbO1oty
HtA4/2jwwB52eJhr2VdJHbYk/1JCe347exUtAa/voMPFnPI/mws7IUkpCaRumnwNo3XOCmfdqOpC
lFVMjQdelwNJpK3ayrjAmZay/2MUQu6iTYgR+wZdim4gUszIEN2q2Ua7O9ELXwI/7/97LAn1qhI2
7mxa1fbRxH+6NfqoF9KP0RJGVHdI7eZBj0rtknp5xKDwTux9GdTsWXyceARbaZr6BqVCL5CUo6TH
ZPlrwuoer/uc7phSAheOunHTSHwKh9YNPZZVxiYKyn3OZ0Wf6Whj6yFOxpzxTzJheUZ7HzJc/LW6
IS0Or+ANksnAW66BEmPxSh7Qz3j6Sltuq9KSNNf7XDszbY4ZBlenv8U4D6h5AZskQJeJ6dAHEXYj
XeoAT1Mzu+ic9801Xm3lCMJLB3NwbHzERTVnz8GtSMCMviauE6Hb0wRu54LhKuvSaXoiIHO7+Rk3
lnEnhJ5wAaPlAsaS9QjODn4qoc2svfUF8t5SLIrjfTUYUbdSTw+j6GsmMIy54DaBJ0CiQV3ak9p8
duDUfDhUpGTytTBPlH8P0uoqwoavkDGzvN/DLplT8q9EGjVqw6/yS0JzPcNgwVYD+HLBp9c+QLv8
+RVnl/Qyipe8dfiWG1/HS30XYevFCdSCpNYHsLD5oR8QgjAAy4gWIsgcnZZHtlpDLFBCui5wlGXR
MBayHxGZTEuVu7pfRbHeVj2jn7033CSms0gu+vHneUCURReaB1QZqQQRWvHkMt+KN5daOkoJO6et
VStbOmXUln8GU2XGFZ8+OdWl9M6x4Zef09LmjrUF6TWcHPLnGTW4/KD7GxCTCskCko2Sa+p00PQY
jPMBmM/LA5eITq8p0ZraIt+qmes2B8b1++eT6qNxbf7giqCnpeErTNy7QlrshCSW2nv1OQGJ1wV5
T5zN8Qjovq1cXuDVYXu6SDxa4qs75Nq9F2ukIz7/Kd8nRM1OEvITeWvDI9khpqtTKejnSHyU8pDq
TfiLZM1e/X1wdlFPTR9pKvvivHpmKv1qebuUPWXF68Ud+V64tH5HRHvgSJ0BVm6vBMCEfdjgPXAC
h0sVikkDGAxjxEgQc45aQdnvE6yVMXRdDgaxX2TbS8vYSoQzMrWOm+HGvFPGAU1zIcWGhSVZtdr8
EdkH1GaNvyr7+zp0y7RVvXMxLDgprsBmi/e+zrDQxsErgaWyXCCYPXO8RzV1r+Wr5jdV5siCHckf
rGZacFb72uDHhL6B8apIdk3PTA5ocOqRNpCsyizA+ao+iacJgapkvl1mHRUySwFcVotQyFoCgJ7i
sXcTKrBKZnYcu2NmTTjSs91IxBTHx2n/c3JiU8uuxeU1/69vFMDqKw2jLyZ+so5fdlfDFdMStE+3
InnUmYmeCwGcxnyQNqK3l455QncCBkueqlcM5dc3fDsWA8nYAUGZKrFwFKXclHbUugvM1nCm3YSU
lHdZCXMnkLG6zaJ888ngXS2JqYq9+BWdgePOqGJxnrAenJs5QpZz00tXLGmLvGewNdusx9O4J8Sj
Z27beghWdpgy7MuBbloFbgGRNHIleoe5vRFKcNexSE5xo9e1ezE6KcCR4STdWCqK8mXm+TaBuYrS
SqcJ82lxAPIAwma7swJcaEcKTmZif6C/oTs/D+EXvdLxyDqgK8ttcBZoV1q9gkGbER1pvNoUzUhW
r7lAZf4X3gCe2WOo5f9pbR4C/ReEbYDEH63KE48SkKhFoQZblfRN14cHfNVdflrYS7hdUstr1+pD
P4VbfkLBIBZ/STfLwnNwkkNuP9fA6JIRA+rTvYERFOuRao7aa/itXETgZ6O+3iZbzXA9xR8QKqbF
BWDGCg/bjhMv7KHMKVpTrzqphO1Onmi1LgcEAgu+zIPq8BqJuqBAO3M/5128AbmVtkFmopSNm7wI
KOGZdpkxhH/oCWx5M2l3QENHA/xz8oDX6OKWi3fap0ouPLdToVVNbBwjbd7y/KRd0uq+Cayb8YeF
eoN4SME/NbU2Kc+l29YTI855GjG5pXyUwx7BSDlzYVBeBoDhzEp/R34c6Kpr7v39jBpXX8Gp9TRH
DwLVa21/c2CvbJUQ87vyPHtPEffzwMmJYKBvAMMbJJCy7WmOJraR3xIlQArz4mkYs946yIjDweUr
/s1+hd4dnAyGMkcAhHI9VX0l8P0Nxau9qvOZk5BiKyarszAUUOameMQee6gitIktoUOxPGBn1MyC
GOSf/b1IE6RfPJ4Kx7zXGtx/BTFeBHMDyDJhM2gJI9mmiycXboohP3umQH3wfp6GPCK1Y43M5YBd
g3MKi+c4q5aHrQ4oY0noIBH1ccXtsab9NnFWm8/pKI6K8aic5llVolK+Qvh+cllfkFqUX5yyEOFr
/MRLS/oO8SEQIZSN27YHn+2vaDF6hM+o1sSLpTTm79l6jj4wXzBfNFY1qJJ14tcQXVUdbVquY35f
6NlShmFVxhPC3sCB7GSpMscysJUjnvDKnwGsA50b1wCpPDDaLxfByD6qYVNBWAzRLt2mYoMtUgnz
W7PwvnaZ54OZz9yc87FBpQU9qT7ajvrdyNsYI5gYzNkMxYF5hD08VTo1ZES1xBB1pZcKIgnWJgbG
cSLlT1xhNoa00Dr2YkjsXODEGD1KvbXffcY4rfJOX3QptYvLqqdzuqpRppRinDANro0CEfaQuwYJ
lp5dHgpcFTNgDGrJHGjZefgwgSEDLBOYJO8qBWfhbWxe9bMSeDb3e6Lm5Thxx0Ou/iRb9ihXayVN
8dd6I+HUehumDtb/asF4kTedfD8bkj470yYI8pAF2iO9gooFCH01Ehdb01Sc2790zfYqBOoHlNAz
PUeSaKHphF7z5N5QoyRmITRwJGdEAi+8x01tiSwf8hTu08K/kxOK9rUj3+P0uu9a3zQXMBjb5m9P
r47XwtsYXBSmPsvjH0lPUQP6ee1vru4nC9Yf4uSTH9eQ2/x47tWi8URTJ37yaqlwNn2wrI3Wsr97
sa1rCq0zAOxroB40bRxudYa/tqGMB+SR/2kWXP104a+Ne5LNBky4/HD22gNwKPNTT2865+nkdc2C
pfIJCJAkEH8taNE5aUG9/QtEGkQb7EuFBZsFd/HK5ggOb1jOlRs9qbrOjsdT76BQPeNBbCmNmSXf
/EZJ4sR0TsdmchJVSvVXJ8ohFoHYcit5HofzwC6lcNm5t7O9XUGhi52mePDuW+iO4xidY5iVxsmF
fz+E4TYmnox6G815WbcMbTFmBiwO7j5bFGJ7xKvvBta3teUoo0mtFQTdhXsCi79weDKs+LKfyCZu
/C6T0BTHUMWkt/Vy4Ub14vxjOA5hDJGpQyyirtpSjPbENdmS+oQZ71dmal/JB+CNI1xlvtfvFuwM
qk+T3Ko9JKCIW3xDmLIAkIT4UXC+SkfnzkIxBG5Nantta2Ky5X3LYhO85tj0YJh6SKPh0zxf9EXT
tKCTV5tAsbCo4eIdzxvL98plnlvtz9IVlsKi61QRmoNiqLgKJ24ZQEFZ5WrmKHzKGVy/KC0xgULG
RXBQ6HjfDFvMqu5Pyi3P4KT88LWs/ITjfZMk9RPxsN50+3qgmK6sw/1fGt4/LtGTTai28dbNHXoq
BS8egPtH22G0NDw5QJWPR0q28YYdYCmsrfgLgmy066ED/b6FoNLj5+6XSCdlXKxbqxUdrV+B9ytC
UXYl3uEV4K5Anx0YjMDagmYpWI9v0Syo6/uTovsrMVf3LxifrWYdbvQAhuiaHt/54onxYn9ylXQV
EEDy+7WNzmbuDTHQRFMqtOkaJ9thC1Oo40V3CrnCe4iDShsTk59m2Ud8NIWLCWQUx62SSNy6lPhg
RrXT745zzToa68yjETNSehmBgpwb+CFwTeQc/CrAJ8X4uJE9hXJsPHELpxAqh5cJgXcwNVy29/EE
K14kmtXlK2M1+MIvhlKOXqtZntJESr9VQDU03HrYJFVvcL45qFa8B5UTDXza/i1NC609VfSdGKdp
8siFUErkRyaKcQNIROcvCZo9wN0AXHn0rb4rBDQNlWBQx1g66ScPRPeL1Im+HFL2z5ImShVnM58n
cIWQrc+DYyIb4iu9DF2V91mFXFTiO84zv+zzryuUGt2DctPBZw0RzKoQx1aA594YDoJTv0vrROuz
dYYnCoHSlmELcL7jcKNMYIZ/eD02WfLPeJZD2DDyFDZtCoxYM1Iw3hlDVBk27OJidZjoWqT6Vaww
6ZrjbJ1mvouOaDKLZ59/aliFjbatklXGSdP0ceAkNEIGLZdyvZ6iCPwNsNDYKvTHFLWctUuPLfoT
Tqx73pn1lO8jciZu8QTOYO/XFYa6LvfAnjKFsc2eBVshWL+eNf0VDZ0jueXY7fgs18vBxuVvh/2P
QZD8g/goNzJ2mDJHHnZKO/tUrC+8K7rxjlZbdp0vM/QpmjrLnMOGxLPtkRBi65q/AUYPNVwNttC6
Dq4fV9vj7lOV12Vc3xUahmAxgwdJr25tn/eUKCue+y8zJggouB/HMAsMS63hFPwG2tTbT0dfoMsv
eASI77zMlH0Sf9QrVk5NKCQzjOJQAsSAO0TmHWdOesc5KLe8K1flJMH7Fof74+JAMr6y4i/x/vVe
LWUoZH1GrVkEcW7jf9BTMPq/RcSJVFThoAFfek5iYuTOtNuf6j4hFzyBClOEeSfVbMlU1t/XYyGx
jM2qTGgTduPDw79WUDwEATQ2RY2ktxLPVdBdcieGFQFH/MAh6eosAw/vBgcTZzt1tGjTaMYYFmZh
sruR5EXu3maXZnsc66+FQp+mOOVW5ZMOmkXtCxmr3DPzsLS97/ihGLD8OuE/X8cfIQ2vEM03JF/Z
E32jel51qNSB4Ef0a91N4Fwmgth3eyb1piWIRQDoKfviSl+iA2Pf2SUaiqeoijJXs6xmb5GMAD0S
QR+90x7/RyZob2S1f+HwGSTBlnCfXUnT2nEsWk7aODgvIXawEHXi7KfA2qpSrBbUX75MECMTpUeJ
zp9FU3AVS3AeHtkBP/zE3Bz0ynDMFx2aC3t78oki7l1Vlk7N0rJ8TS69cbAMkWDkwTApDVJ80K9e
z09NT9D2UrkpAhS2KAwKxzVC4yJtLjRWtenF0TjrvSynfW+XrMyRVlOSkEs4o+vBBFMGNM1vGhRv
/0yBKaUUUbfsDa/zr/RIYjffzLu2uzSxAMNDyV71I0dR5w+2aytXYMlgvfeSPi+Iy+xzP32swWRJ
fLv03j9Gf2TnXGtGDYvkgcw/f6LySPI+LGoFwShryJnsjqbtysq9mRVW0s+4r5MqHKLQhdDPe3lO
27XtpvULVCU/WxS4q6RRQh2J2inOHz9Bvk7GvK7TTx5hjydaGSKGDisvBRt1r8k9i0uG/M0yb0dT
8lfcBzoepsjDeCn0ess/U1Tzpy1heGnAWYGUb1kgSJ4gb3lN/QzEtAH39jBN2KVLNDA3atCU+PtU
1qx79HC9YkUR0IiVhLIUK6SU0vhKfcoVkFRoZI9CE1UsD1dpBzGDU3djiDpYE53likqMkb2RKYRQ
lSfMWk1tYd/IaOaLUhhTX1BmMtkgPSpLxD43cbetMcXxxl7tmJaC/dkUVEbpWuTAdb7YkJbJctjn
QfwSw0gGpxNty7IXJ958tBmUIzwOoOADX42HwLkJO+diVR2DTWO49UIZWcuvAIt1m9GetyasFEg9
JClIOTegKXlM1pNVZxfYGDDhXQJo4CQs97bL4f2c1byHrF1RN6OFOTU4m2+2GW6BJ9TrkDBloGd8
yXfYZD2oFw1QiBQ8nFzrDVyGxOW7HxSKcPR82UcHI2BwPwDNM+gTjwSBWm9Xt1nbB8AwbmDiU/Ba
sbhjXR+Y+P1mWrlhkG9HDqUcskqbPNKu2QrHT9i7C+Il8S+q8Dxuy6ERsskJHOW0MYAUbFdNQtyY
TfH9yfxqfbNRfOL7DdSmoZWs1eTdmTIoIUqfuYqgf5pt8OHdgoi790u85YQqCgaC07AvoeQjjvlt
ldrEsqZkdlutIzTlUMlIJ6IeMLsvH7xOY0+nZT4RkRr9al5EszY+qp118AeoqouaxseI2NS72FWp
IUPbIQB5gMm5PcH9tKHI/JjcSpj04xbPaEaNZrkYqCKeIAC+MUDiu6i0kfYr7TOa6SroQ5EUeiVA
persL82uIzzSZWrcRYQ2/Ke6GP+SWYDfsODBV7BuDHi3svt1FOUnf/oN+l6YRy793W/FhWVVCH70
q+u4LBKTYvuwsDcYxCHS6ezKPFYRjaVsKFaTUnUBEY6QZ0Z9+w0tHD/8qrUdne1eQG5OTdhq+lRP
gFBzdEyXNw4A41g6X8ANyhxLuYV1Z/c822P2AiwwkWNqrRN77/VAtGBAog8u+gYfBpBkB7iisCfi
6jr9rTwKyD/+rYcvFV+wLAnn3BrjLXhiWdWtNdL++6q/L1HWdxWpNeix5EhaOnxF5RzIMUhzhfyY
68UDB1k0z1klI7VMGbcjqEvQ5nVScw6ktdkMlLdP4/hEIewuEDW3MB63inKflc5N98de+g982U/N
YsRuNGpTyeTQPWrln3k3b+dBU7+lsAOeZIFWyIk+qjN+UQt5dIdPcmEVxyN8W41PgfyqYKEewkO8
sjBC9d8bbdoRvBZVorp8bJX5OdNAAhnpbIFYt4uVX4uE+d1SLTyL+L6xOKrywCKzK5QUVcpbGAdD
hvCizhQFivh+KQOzVJlLdoqP3AzCR8LCpKIQtwW4cejybPQj9SCx05oTMwJeCvYxLK58FjhDhGl7
+EkFlatpu8TQ+rUvqr69a79wab4UIRAgXpugGfMaOVA+JPwQqCCVePFpqs/MM6OjABcJtsEGxe72
ad/fPDF1GWxFOyHDms4/U9BzZ0zsGigOWdusv7fP/N04iK2u144dLB1bcqatoEvPg8ucwuPphJOh
LkGhQyfaDQmz/QnoJMjps0bdKcaXekrKx7IzlDp9mnpqVbnaKMTH0tinjkSJcyLG3jkqhjy1vgrQ
0FhRm6S21M0C5OwypRzQKCvxCgwX6ELbUUkiiPzVZf43zO/iZSOHxtaheNSVXeoLz3oF+fNBTadH
i8C8JA5+kAbNRAqFZTLR73/PCAQ3JW8jsG9itft+gXv3vuZ+nWvdS1O2h3QqkuSkgy4P/YgksbyL
vwAiSresL66EPjrzQmJE0pdRSQpT2g17hcFNQTOa9j1OnkoHmgntzZkuNtAVsRR5IIUYd6xLzFfA
8aWiAbuE/7UyT+NNMb3eNrbAa6dY75vauCUf0uLV3QRkIu6iMJ9y0KFqrOhmhhbrsjaVhewJyPQb
TaKI4KNXvfX0iRIJ1MMLK62judq7gReuIypjsumsaTZSW6SL6e/1eQnoEwS/Aj6bIDzJK7+sFuUQ
xuwbjdfYK05vg60iW34/Pyeqfs+iB2fxhYorR6B5ogLRiZ2irdpXg6MdkNG5pPX6GLYg69qophJR
buh5yEOEjS/7akab6DI6frtdIXsi/bf7LFDk7X3GEWNMLbqrX1sDXJuMk5lCjvXc5fHp7RXgct3Y
THxwwLZkkfg8W5EIvslqrmIkPMoA6c88jSJNxUy0WhTurXlSgJb9do9iMJNk4d+ElA21E6Q1GXb+
Spjqjkj9Pjw7HSQV9g80o+0f0sDwkAAqi1dzfwHsAzh1xKWg5CCbuamDvtBeYHCvMlsrcW0q8mOg
mKczMOL1HFGdh19ZOC/0Le79C5uFC//RbyaTGAtOzGNKCZja+v7bLyt4bY513zO8XM8JHq+6ouYL
Phqabx8WaDhMCtWGNfxQLy1IDwp5DPi23GakitXkNPqNiBaf5z8uttLkqzZPP47qdGqhQP8JNwI2
XG3cVMtHxo4drlC0TdCtSzOJt3wsaysahzXNMe7nu2smAm28bm2fBdReH5dZcNCX+D1Gco3kW9FP
zWUukBiPtv+zG+LiIKBJzH4PLXcfdtxuQWLcviGtFQ+NvfG4FnINMmxuCiYywgaZJ9BU9O3I2fEW
xqjL7zzdwTrcr5HcWxZXLe3Ri9l7+E+tLIIBuRMX2vQ/z/vhRm6+Yr6CSVTPtoq7/rhrJpfmfUWo
EhO22c9Cat62LjZiG+an00m1EzGPv/nTH1MXit/v95haUypIErEiPzEh/NL9M5PBLwI0VUsuydWO
65PcTwwQT5Xx6nfyGa1EBBScpvHnRcnHznMvTrzUAU7zBae0pCpOgdB8v85B3URpI9N22id5HYFS
PF84LikLyqW+YiZh1BFx6FuZgcPS++8ZiaYhl2kfx+IJuPAMDfJHUTQx+vL6DdrrIdYWSCFnaXEV
zBBa8fSL8tdWwm+mZHDwIRJyL5FZwEXRcxh6fqlOqdArLsvXVKnsdEfberiT+2RIzIiDoo6+HMoA
Toqqsd8JWbux2ieVu7/+MqiSI+yHoCLoKmQtivZTUaK701RHRXIzdH0+z3qvCWuDfc3F5dzjY62D
bA6yHbVWhVhGgI+sVFrfVwOWqACSFrfcMuN0bZ2wmt1qWG2lHskz9t1xXrbsDElT0wq73roDGtX7
oNEJdsNsZq1ypeoWsApTaWAMhnI2s+DYghyH50VS3KgvaJSIuvTqp1AWj65addkvl6OrAlx8pphP
aHt+m7mSN8yFSaaL/IbXSDrqiSIeRbAIkX9hwHVY2o1MCYzyT6VJ07ScJQHGLu+8rXDJUqs4xRpw
HZiT5IOa5mV2JQOeZdDkYyIU4YTaoKzrnLloOMnBjnoN3ZVVEfypaSYwL+DyI7yL6LnLMTapaBYo
RYhDqfYRHi9N8IDI/FJHgKGml6nXov9Tkfny9gg3lAzztJMA336IqZ/UYiIJH91faggNae5R8X/D
1zKIs1vM6wIBDr1ofa7XVYevNkyMSsRP1YKKSupejNifuJx4u92B2cXi8YnJ5CFS8CuO9q7km+h7
qvu5lvObHp4Qt24tbLErgKXGXCD7H1LvzBnk78GXF0rr9T9Z8647Xy9NHFFTZLTlDp2hh5xQWfzE
4gIkbEvSnbBo/njYID5LWp/7NzJxoM8FA1odBrN8KT3vg6iVsltKu5uOn4ydBWqPulptL8KaBazZ
rZ55iSFOvrqLnilK0dhQTDFjN5IBgydcX+dHAqpiXslkuHLCRrBXT7dhVW9R3P84YYVuJnFeu40w
azrUnLv7EG1FSL1yHDsvVJHonPLtzIEC/FO1lrhdE+ZR2oK8qsV7ShWtDF1bP2fUbir7YBIY4e4T
KIBWKvWoT3aoXfiQkuT1W7HxhnZwPJ7VVIpNuoN1UEfb5D2sb2JI5yHHVkIMBW8aS7QhZN6IA+eo
h05RieXi0wKvD2wkBiEFVd2pd/VDBH4mI0RSglzGzTGAXn/ZqnmK2tur+Z15+xJ46BV/boYH5i0K
/te6nD5Klr8/lpjBXxoYJxDMGoJVXfNeswdHDxr7MBc4cbv0eolM/Wd7M/YoR+2l5Cda/VpC/TZc
Bzk5Xf9UIHFkzqxR4zgy8lM82iycltezxYuxUzrmbRpumai9HzfIiLDqUX1wDdIQfimMYh4dvfaL
qQxtN9u/4oYuj4gzAt2Iqp+Fh53Ra9R90mi7kxR41vnGACPoOhbV425zP32J++IYCS4y4OxQsT+0
rveGU0/8XDQ/3KG0vBY6xZOZ32ocXAhpaFaMsTh2a4g8J1Lm8x/0B27OVikVTuidY5PgFaToCWmx
5UNp2XGivj9oosQN+fYSePR7xph26TiztHL9giw+7X2OYD50tyjA7SHZ2wXPtrr226akK0m9h0YE
tZ7AIe/5h2atoUwHelxgOz2A1mFF+RvC9IHqFYtrroeuIsU7zOM9c5CRoC29rjTfyNTZR21wfvBo
JD8Iw95YQJu1CNCzHX7EDAPUb9dIhkG0K9+1+YW1CPCfGv+c7zeh4XBQnKGhlri6G9YIOpO34KnL
BeZbelWK1AbBuRm8IRT7dUiUpV0zSz0S5ZDyIPEzMd4S++/IXCJmzZuYPXJSanh5si55+9Ml0l/t
YQ3Nl2t3zhwdX3ML4HH4u2Nc6T06rGdsw4+jxyEk/h6f/GBHq/9wXm/voM7m21SjKn+ewZAvCVD3
Dd+CXaxsUdJTQjGHT0DSul6Tqy4KIGVyeglZC7qVtgLm6K+DiUNtxSaliwLZ2K1VbKWkiXzYb0TK
w1xLmvvpXlxKqNS6bVY3RPBqJqSUwMhv29SaCHYMsNyMEPh9P2yneCu01wOAYQkdn9MOlzdlg5yW
D/VOD+1AVXbysask3kcIDwVYHTxR6t+fJBbSGOyvYnLS/4rc2kISiZvv1q+m571jwkbn2jgRs6p5
yIWfETC1gJ+uuEPFrvaO4Pj2vxUft790NODnaWnql+hZOKY6JRPFFW2ek1diCpiBqiijKfmsFbPl
Dt98Oy1g7X9za2Ya46hN1ghifT+NC2dE9jjRi65HZaqIxZjdULNm7go7Uj8rBP5FKWekJg1trvj/
aPjc/kikzhJfEMobgI50pVDfJ0i3pRTzMmgkwraYtp+I5ej/x5p+RiiLTAapigkvw+sXrhgk+VLH
hJtDT4mp8ogxywmdMRlrHZik3HosqW9uh3iQ6T+BvcJlo5VoOBjnrt13K6bbcpzgm+IcXwUEu+yd
7pz74D+39wtJM1wE0bBDp+7/A0aC9FSosHHyzgi0uINoOzXZUM3ii7apWV8/jwI03mP8W5zbEal0
tKqgoM+SfDc3gXpmheOkuerfGHZyrjdI2/MRf+94FYLJbiA2tmcGMDmvl4+DMClgelDjNfE2fKIS
v666tEjcFcvwP2EJTbRF09J+wpsbHHS2RF/lQHqh9BeY80pKYDZCPbe5264GzOuOqgv97o4LUola
XXMYXpMfN3JdfYVtHkwCiKZEzmbAOSgIZX7W5NcrSTRXjyU6dIdyykHDfIf1qjR+WT7LhuJ/izJT
N1+Tm85UwbichkISTbv6QY91wK9YcNGEwXwq3S1gEDXhCiiBwXdybxGN2IcHfqR5XKGsJtIOff3o
gkxpjM6+V/aTL921N9B/wFXzA0jGhwZFl2fWvhg4JmoU1PH5NdMv8xcFPuBziNpXLknNLK4Gk4WX
I6hSbUlJ839PwqYg26gmTtbN3oD2MtdrfsQOBuLcKQSgqHmMJqqHIM5B4nXh3CNI27lJqjdcqehr
7HPK1LN6AJ3DaR0ylE6hLQY90F9gHdDb64H4MQ9JVcH+JtTQhTjUymsWgPk6bqFvDK5za/TgDnYh
Y2tvGyKpsPYdDz4p/9vRkUhl+5FtUE36M4UKNnY7j6qkAJlPX70Qgc4lb6neIEL19tXCkfVpOqhQ
YcLeyNnZeE7uAKLY4gfrpwBxXRamfwpaAjPTg/ptLcj4coi+g1EfBHC9ou1SiUx0esl6ojyRcsBU
d65WpC1G46jJMs4zYxkNnx8bRX3f3xrZoFF3geUKOqdvVzadxtQC3iFz9qqOKj0KO0VFHYZH8s6A
LZkkplm7kDvkDE0G5Aqnq4aao1zV91jIfaS+cqoUBp28gRRxY1i+tVXO8KJGB+ZHqw51rjzSAoRe
l2Psdv8N/Bi3sT86Ic1rsIUcz8G3iDjW1jwSbxbfe9vZEe5ZMc43+CZrh4S25D5BzYCCBsolXMDt
7XH8Ic0oIV8PD+wCI/Lws5gNQg+szlYdSF4tQFWVPF1dZfnYnywe7Q28ZNOLhPRTDSd8nnSDlFb4
nyjRrQCcgac5FO3fbm4q/a7xx4TBMnYbNy03EJfveOBI6LfiOC30eIxJ34+MvQy7bIJ9zulXUxog
Kb9WA1CNzz+rnwd7fkxXTmUvE6isr8PY2xkNBEWyU3j1AVefasJlyFNoxjrxbKU6j6LNfJ9KThEy
XeMXOrbuwhapVm6bR2J8wt7PExQbUok2y+up1j9M9uUmxPxtjn+v3zTV1T1iN3IKbnzpz2vANgHJ
MJjF2lvIabOPGGGQWtACn3zndAMFqtkO2D8Rli5w+FfgNxaXJrsBZUDWMANaFDrDtkKlGWfnoOh7
g8OyhfQZUshWMPMU1pbx9acbSvkt3LhWtoi9S1rgKlvmeonDyEaCSQgJblhv4MfTiCztldmkJi7u
9zqDaEQFmn61dPrF+ffdsB143zYceOMrAAPcw4hNH17l2Nh/HS2tS5KsxWBFHeKgNBdr5pKOetkP
EHPfDqvwSz3lNClvoIZkxtnfb1FmkBTV11P6ET0LFiQKyNYJKH4Eh9sINz408ZjYokk2/Wc3cme2
j4zOcW/FbISEH2sk1lm3kXWnJyL4+k/+74E4z4tDlinXkc0BmIWMg/xtAzIAGqiUcXpq6XjFvSGj
DdGEgfIeC232iZybt0pRbg0ifXp1jTLWTehr6tLYyebm+lJXvPbfYVFXa+NaTWqUZaHwjuHo1Pzc
c8kDO2bzXwgmhfCok/RE8NqvAYv+feRGr2aTVdTCEx+3dSoUMLClA4O7ImhGovPGoTRaz31BSVYu
6Z4cqNFtsWxiBljRdo79x1qMSgm/L2aiqe8VzbSGJPmqougs6iXKxjtz3VDwdyOGiXPD1Vi+DAQ6
T2fKJPut5ixhjpvcRRgmu0+0rMMqXq+PBAcF2ZhIqidBp0cl32Ws0ltWyq7VnDaj9E4sIBfES8XW
g4ew3Gx/+UdJPpOJMKtkz6G47zMQn+OMpn4tiNEx2DVepZRkDk4rhgr2UWicrKW+NekvGRG1lZWn
E1+ryIyh0+6zgsHomstCwD58JI93hdhQGIjV5SG2CuNAKsKJohZg77b0RmHwnDTQ2QzFeezEEvQs
BnheB1H/dgFPTtxMjwMLwyNYcw95mhiOBB1rN2u6xMoeIYr1iCsmXEaSWOFcrTNjoHzf+rYcQGh6
z3U396xEnjgZYuDHRjNfHO73GrkrvHf46N6aNUv56aoLNfGDPPfItiLd1TgPlulOPpow9I8tlk9h
+W/EdsDzMXhaUr9heysl1fgausYVMuMDxOnH/ohyfrJXililQgsu2y7QxjcJzwowzmgEhaqY9dwi
oFFYyNh2+kwzqSsWf1iX0kwJM2QdJYIkH8gYsuEOsC9vRceMDE4Peh6B2J/Y/SoXxPXVelsxgizy
0mHVw2a1HJFRFCwWqTsb5+GTcGwJxZ/LyFrPaLMAD3OzuPk8oNlPx1OVVLz6KfAhlgDt7sqdY6Cz
Zc3ayy/rB+w5aIv1kgUde3gWLlSzED9Mm5F/sbI7ijuuGvfEOWvjb0AuhIFsyjjwznsvIINWy3oH
8SIECOlK8SkhXxTMUp6cSRtICAodlZuWiSsJJkq8YaMsRkOLTKF4bx7y3kW/bbVC/O1PfBdNQRoq
g8x1S/cCwMJj9bFpfIrklvhJucxEx14wuzgdWOuOhu0kTOA/c+NmgWR2MCuXA8biOZ6WSShYJME4
DhEd9vdzExcLne6xKOBWtqQ4LavEIABPuuzD0N5zWj4mSZMyFXjt5lQ99ni/Zb4PKa22f+u9jB2K
PvvMifBob+KBKZxDcHXLOIiHyIt+6O2oKTyPjMrZWj716QXMdnyQmwxzAFv9NlbWA71ZcZMUMeKW
n8rGQV1Xbnh0t8N/c5zKypgyFzgNkRFzs6dTCulbGmD+Jqmzh/HrXpPSEJPfvgHJF8jtTIVhDonz
nDV/C3DV+Rc1+iABGrmsDKbKN2B9DnSH/HFxYFn0qKU7IL8HBJCH7VdbYJ9EYoX4iSezZ/OEkuOc
cSITLJj/h2HL2+mhA+SDDWcPlDUvKs8dCH1+EnQJi3BwOMt6aUeHiG+G3GKN6zbTE0/R23Y+FW3I
LopA7W0D7vWiQO9BS2q9wZHXglmlHKC22g+CDgJJW09CRxU3V6MJ3z+gTYl/O4eqBUiqf3AluZ7c
zFPPKrFy9Io4Txc5vaTUsy4WvlZrV7ow5SldcdQTXmUFYJ6XpKDqNAxbG+gbRlctB5GJYl81SBEF
+X+vqKZj3+HRjhnznhjb5iDhVy8u12VMIDZ70Tuq7n8tLmN5acHunrnZmJDmVbPULBiEpGQ21N8+
5q+LEvh6Kle5I/9hymYg4DU1YZvXKx5qZPDnegjAyZtyJd+Rd3lvU8fv4nqg6vt/scsbZwECIgFH
2aGb8DbcI4LVK+Xu6jmJis9ncWhQN3/2G6P06OsRnNl+JL3ZnS1XjH3mNybIjiagbPPMChgf+7rp
iyYO85cWxQN5Cgfs/s9Mo6RmEYSEggVGMfq8w+/neksSQ5a/ow78zS4mL7Ejva6o03ETT28Hzwbn
nZ+xQUp0UVY5L2NckxvxLkadoQd3Sik9FhAHt0nty5IhkALJKB41QaSai+2SRaMadp3YOmLJDgJs
iHI7Lz6YydR3Re2nZtlXcMZvwDTM6TkYegHJXRFw+WDOwHS7kLSZLnn6rD7BGSKyjl8g4PJwC/ek
0FjcPF8IApemszc+8HTXFkwMIxkIXSiexPjLxz8vaKRTeWHiBgFm6dJ8wjhtIJT/bjnY9nhA3ZXN
2kYsNAVhShfEp56to2bJGhM9mQagKZ68J0lRTJryi2cHUGoXC3MyD8oT3C9mW9HhkvWpD/RYdUtt
8mIPVpZm3p2FqPZgE+dhZ2vQ03PpTX5oBukGzYpp56Xe2knoKCiTCJUpSMBIxbr7X5PKiPFRyuMh
MAC/Q4kEOb2sLRwC4HUPm2ipVD3+MB8QP90tYoHIANS7fu3l6dMZUXb7ZkbyX/g65j3o9DcRobcj
LmQloNnD5mS8Y6xP7onjQFTX7+F8RTWTmHGhMewLfR2Dot/BNhfGV55+AXB3zvUF41OmumhRbxUY
UgvnSRTnyjcFjyXvwvbxGY+NCgHvxTS4nt3jafdWuLTagja0yihpNMg/hTt8qz+pRDATGKlMdMoK
v+tvZLk8Q26QpaShyd1fDTo7aG+5H+TqhRSQNL1chl/F/ATM4QRTtC0ASlrTTcbCDyJYvBevEBbE
ESN2rCDkCUC4Q9bSlCwMU95DoIxGsvkgGw2aBkyHKwkKa7V5mGi8mrm1pdg+nHyqO096FN1GoH7n
R1WMW6dNc3vTAYxLUHHxB439YaRy7cShvJSv/4zF8Rhvab8JUKe9SMtx4RiGn7sFPZHazKJ+fOO/
+zB7QiQJXmQv7XhrVA+u9hBPPA2yRmVGTFb/IH8UZGf53CAdr9mfJYpCHT1mpLxDrZIwnuv7IIpM
k3Zi9ox/mQnuM0X/MHzMVLLGmMivc9FTC5ZIXLrJwMFExzCaCSX1zq4uAQO1HQH0htPbcVDqMmk9
xeykrLIwEjMGGPukCXNUL4DxcVVO7To4TLCuYjU0fABn79eC3jyb9/PCWfCzd+gMmO4lWwnCq5D8
vNPuJdOKZDluAfKFKc5NBb0gyXh/26cbQ2ToeHNeFQbPsYEl1tE5cDMyVPCKdAbDE1U4z0Pr103R
dDx1lcSCxEWtdSVA+Mm14/tugyrQXojaneX4Dtrz3S9eCUDVdSa5JtwlqS9ojjDU/oHFQ9Q3PCR2
b+XzInla44iR3s2In2czsdpwhrKvCpiID1wWruj0rVAaw4ZhtBWLz0jK3p38/wqiIguSmIwT1l6I
IncflTuiOwDdm+hJ6RJLX43hsFmL7FFQOqPzKXM/8gp2Y4hIDmB/Hz4kW6l7MRkrh7UAVG09zAFq
JFBz+XctNLs7rqk7nC73pKyeLx8WQKN94cHDs2GxhEU+sEnrnF/b32UTmi0aRB7CZ6hAo7o/CdmV
p0MnDra0TeAv0OeGpSZbFXjiZHykYaAGe+DJh8G1Um5pSBfd1rGZtucLhLjfj6kCKCAWTTRiJTK4
cRhmWQWlSUrMTbjg33aYDzpGFeguNM2oQbS41u5JfyRX+ZfS70394LypANrZtQSroie72KSgWfsu
ekCeMhEIzweppnvdKnuaCLcdH7ragiyuJq8IF2fKjPnLQQjyjUC0r2tnNP31ajxYHYoIa+HCq/M1
SElQhueMXfziZ6mYbQoXw9Sxnp4kbB/Chjn2fXa9CuVkAg/HH34U+3HKZ9voEo6ONce4kE6DOH7w
P6YPXlDtEjnClZKrpAOrqBBBALYLJaIA7h/Thkv1Nm1EfuSXFCb5diFvqrewEohXtt/Mgm1ehGsO
f4eu45rzTDf9xPWkfPDJJE5qbY4NvQERwazdH7tjazw4X+pAcfQ3Vovsth3/gU6olat3ApDbkOp1
k+l/ltha+fJDr2dqqaVFgKBGl0gy0kgzdTfJ7cELUdKeHnB9doDsGhshss7BLWusj3U9kvKnl/bO
VmqU+BeZ8XWoZYGoiTgC3pQuPrDVpu0/edJ9MAL99t8hDKJ6Slb6reczLQD3F0rHLWCH60IxCu85
zTjl5Z8DMZmmwPcrAGA8FZXHpZclYs02kl3uHSuwwi7oBFfq+hMl5j9g0hoNuM1QdGRWvHiw8rmE
Liv8EYwDytvlWCY841N0Fg2ClR+XocAb83c6q/e4H5UKtARzGCQ+Fvf90Urew0/XV2qJ0vRKh0+o
VebAlLSbwG7Po7ItInH2hmBmAHMVkbYMMRTRCpgCd97Ex/Wt8aAL4Kc+eAya32QwjlMDfVQ3AvwR
Xwnrk7xrNTIB/cUmvAUm+yllVUnAW+X55O6gCWik46iOdaQ7aFksSWhiJYG9LV5VbPFeTxR1w8Wk
FQqXDRPMWQ8ImxQsfBOBqGi11E12Q2ip59FHmklwBwatrHhtvOLahAcMZd3PNSrOFooTvAUFzbbr
0ZyOboZoEvUlEReSycJR2MAjpS1A4Mf46esTCFvSVi0MJsmtmzr3Gur+cHcPgjnRjo3Yzp3BowNr
ImwNuqtEyXDNnDGz0BgPeCSLFlPLvy3febfffmYQCSH9TlGF3H927Ox9xlycj+OKWmsUKErLJUi8
zVjR4BpEddvt/u1RrXO1uqSpW/ExqP9mII7xTCwMGMbRUpQlcr8Spv+HuCEBsdZzn2wsTETNQGmH
y95Q349QVt+c7Uzbtrx+NpFdi2Y0ghc12Ki+X0/dgegFt8qeC65qmjSdWxLWmGSqA8RsUfzhGbmg
qgrdP1e/BsC3Yc8gcPxuFsqDHAqSeMzBVcgiZGx+TG4yZuT2zl/qhrj01Ew5LZJzBToitqjBiAdG
Io3osn9fyRCQnLRreejQbj9iUR8/3uOoZ2nrsdEF73Y6ag2mn/Zy+NuSrcQ9AZKOSvIsmIpeEr96
40rsXI6Moq7gRSuAfwWY7qz1nZiDNfeC4XVTIqzAwdmnYmAs34+48Lx0vKGZTjWP4nFi2L0n2jLs
rNCm6FKhsUN0xUbWUDdqZWNz5veqvLWs0MIF0cEvbt+QV9DxL2GdCoIyEeGgvBy1oeOU7q4M/sQZ
65DqEE4LnIyOWZMcmmPJJ5f3jdNZSpCBiy4uk5OzZg+zkBFuiE8ig7TbOiuBEQSG5p89UAjTJvl6
x0ths1upzSWNOybjHnnWvYGXcuDTmMrD4nnB1fFE6pSWuMPuDQOzfVuGklb2Fh4O3tbVlZr/y/kE
iNc4kOP65eu/5qFJE6PdHF6uc6RORDGeRmIdYE8soR/ivEY6eSxt/crMDUifA0VZg8Dh+Uq1Z0n8
8fpxxuLWUf6mGkWKJMD2xywSCCoVt+gpaVg3XZkTw9v1kaEHaKBzYHjXKeYZH7ops3p6hdek1xto
kYwcnlYZpw0rUWtF0V9lcyiJpT5zpjjt2GpAy68Yr17ZZz+4BQsVzo0DqaTRiD+sJrI5k8/YJIwx
rUuhr1SyQ8GwHyCq5XPa4LFjFfYcvFhOwjVZrJUE69AClEtq2FoRB6NVKdmvgxcX7s4S9z9vExRA
vajtxAyUlsfHBmtxk1RN9EtbhXDeAV3OkpSyHQFFOb/7JoOOxetlpN6iPtCXZT5YbAj5x2mxVoDF
ufVGgaJfP72DdUOADrljakNTeA/b6D1eWiM8qN2bZTY0J5S3fkxl020eD9+58lpYs/tlrDqL7nrS
D92CkZ0MedAi5HhTrAPcm6ZFVJJfUmkScyHb+ArsMZBPv66b+Ei5vqGhql4qOPRtmllYdN52rXSq
QaTuLF6vqCHl7RpDU1si7NYNSwaOnrmEIB51ivec+9bIyb+qX7KxEqh8Z7x5L/C0p4OFhAdSviKw
aZRLe4EU6vnhRXoc1ua2TkjJAYKctHLNOmfRHJWCXYbp213HIyW0YJReUdtmkoI7PtoeEEsRHQo4
9h1I0EwqRrgWKtLZBEwgRYREV8vmVjUBo3awn3SX0Svrp3n5PVWYqWUPjfGQwu8liLJ7GBxKeueM
aqGQXuwBLiISCnDPkoG2HfkSNkkMCQ+R5uYJHJGDajN/YOYdycCmCFGrAiZxBwUVaOHUePo66HF9
T3IUCH13NWDrGrpgpit48vIdgXARk1iNAcJ3TXQj+adPRrU04yNdK3sPMwNpw+rP/TPk50SvUP7A
dn3+wsb3gdnBo7n9ER5J5XHoiXp3UOhiLqJOZm0s4qg7vPGCWszpKSsx7IHeUtDHFpbLloGYgy+q
Tc/4tSWnxMB/QMWKjeZfyZZiM4MuQkhTYOP4qwK+VGq7WrTyIT1RotUj4ixf9rA0cP6d263ri8Df
pmLMnZ9j3GOpuFR0SWKAkKrj6n1rSV6XHvIU1MCDyB18xsFjhqoFnphMUuAPslbUrtK/lVnDx8Z9
Z+DB6ndR14Yrh0nmU9p/PsBz6p79MFUFDmJi634+H5IckWFLp9t56M6dbzGrI3zw/onef8Ve2zDu
ASdA5QX7la3fKnLF31W892gHjwcypD8cUDkFrMZEHuZJdtFTN2JoPfXEhqF+fJJVMTSCicNqGGcH
8YeA+Hn1LyH04k5p/8nFDNrsYK4h4z5jBd2zgznlcsi0wPBPnjhhjBdW/4wthyMaLtSyKjYhFG2R
kOVslO88LiSsjw6fbIR01rO/7CU6n3EY2TTLpa/iP7Hp445NM/UG88EuRZv+qmB35e/ATStmLnBG
3dVDe3OLcvGdsKk7Vkj15RpVfl61qXTtIEYftrxHb9qQoBTW/czNL3iHpEtLRzMPhMuQlOeCLizP
sumbLCg6UrMJ0+ePGpuw5l44og4FGI+pb2SE4SXx1ehwwHgF5sXBi6UgvZMT/LPtRNWyu+kEL3m8
08ng+sDxwO3hjpu2TATUqWyRWTf/4macrZXBVXkGc5Co98EHUlSaWDGu5G5BeQdSe+2h6xtww7zb
oPwUjH4dGa33e4WEt8gLVrp8MQaPXh3xYSV2t669BShl4P+1r+xwgroCuzNC2wvFQ9m1LTQBYbkj
sWA5HOA3yC+ByEhP2ffAu8VLjPO5mRYWq6+XTkHkQCUzWJ1N3kxl6pEAlH4CKKA/2R+3p2G4tbOH
cDE4yCC6gt65DOpiIL8X7m3WIv+89XHCbbD27tkTyEdM3zDTEhvTh3lGggYttmohbUhlJBUzZjT+
1A4nDuqoGXXPz21wZh+z52xNjKVXMWW/ogEGE49+n5UT/Hs2AzZIYObPWbevGv+TQkct/KQVLgCs
S6mHd/mvNsRD9azfWIWuDRymk7Q7qHYs8eeHj07oxuE6N14TRjuVpDFX7Li3/wZTXyqOQ8cDgVQc
v1x0a4XulfyZctbpKtiNgC9vrVFJ2dUSG1IhIAiv8IAU5kGl+na3OHFbTDbP8kz/pOvwo602ArW6
rI9JNBnRkzcCcXVAFSp3MYj7PJ/x7z6MRHIndA1FrSO/M2WX4dHT2LUJWS7Al5CzcVYjllcYAFC8
dpPT1weudh9k/Iqn62c5w9V4jqKyWFfzlAw7wDYGjHd62reuNwKGzKKy9K+rhk72h3TDeIIyaQ8p
ouf0Fj5kR4uCUtE61V7JO6MGznq8Saxr+ox3kup7qxojU4ol/MR2K1O1//D1LGeV+boYU/lfm3Um
eCb18h0uietoQeb8jqwl2oNqOtCTHxr4C8aWGkjrFMawzUMyXjmdVtlZHxk50EivuoXIwLmxquXU
EJ3ltd59DqZiC1Db7xCvFfeX1Vo7971aJM/hwGnwP/TYfQi9pvCmwJ9zKn53mqaCAzPOIF2f0OiS
buk2X0G+z2mjllrleiJEAB6oVAEN+Oprjh8+s07mxy2unPbKmmsmtr1FdMKg+8II7j9VEfDLtczu
jreR+eBb4FSTCVYNoQ+bzWDuKezWc61IsDHn+9s4bcK71XKRnb1Mhvskh1AnXEy5pYStL3s8YgOl
Cufe9QpizvP2xVkllMghpGnyVTJcFNUHuzmPngDKJ+pVa33ZGh90H/hGosFYYjMLRdEggv0zYxgU
F6+dHCQOjWGQ3/r+eC/caMIX1Ges7ACiuCLn3MpJxzxAQRqz4iUuuS90nTv9vz7kmfMTi5LZTjjf
G54mSqAC+ho9cq+UqbLSP22kgrZzu+KYJ9j6kzQuhFCzkS7C9QQ6XRXoDBIqwN81Wbbp55YDdwAd
V5YZQs+nNaOnwaJGoAQB44LWpU9fV/oKIvsaszKpA07ufAITJ82KTk8ZbScfsAupiS0RXqRSccvB
IS3xpWGUH3tQpDOcmkODU8XD3A0+PXAGqSVx+xkMZaHLLclG95IhN5eLevVMxhmT63Pd2Ryaaswv
pplRa7t9gpousQenFyBDwG1GEtfsm7+hqIMjTUviYkHTvwxncId6uCnVX3RpXhuTom2OiQ1pspEJ
chH2gonS3psR+ZkJNiRDwL8oEhDhcKXG1GotrSJjdW30OVUTXLHSPi2KXmvBpl6ZSXdiowbueikA
CcTX4O3zY54ojY9wDITv8Y7HTxNgzEIjBwzAGBKQCgjMeAaJRlEYzfmXOsIioU6HAhV1MAbVyYfZ
l3itbqnFTZEZD46t9j74XEQTf4vKcaDTBIYXHk8fCMKkbe8q9yVL1pCHQ/vAAAWPhYEW2ws6VOZm
cNMT7fRJASwTQ00OiR/+vlOW8Fy0B0Z+wQYcDPzu+pcA/cApylubRNEK0pjZWiB+HiMR+msj/PIH
jOiY09uI3Rilkni6KxJLrO/pKVEJHmvkBJIgzgLxLZNID7Fz5MaRUSG0dEDMw/B82U+yMVV27Yfs
uO2M4n9VbODZNC5CyK2BlJ5y50Iqh4LttFNjOeaSIWbv7Pxw8hzyntx5JgqxF+wi7bZhCv2hwlP0
MJAYx158BZb9ZtViEizPTbHJ5kIcrqflYcuCDP4y7ZR8MvJq/f8RL3A86D/L58UcezeU53gL0wCI
RZXbyroaeTwxzJ+HrRVu4CBb65Rx4HhdG5toDGxsdP9SoI8CllRa4wH6WwsS1Btq3UjLC8JsQtOM
DnP2bzfzOQkW6AgiDMEUF+laBfZiWOBV7lPBMTMIvUsUDCrUdStqAtPMrieVyuLCf4hgnuT1iBZR
/zd062N4+ucQbZF6JGYsvD0cXK8D4uBQzr4Inkz27/l0VkHy80FcUu4NpSkFJa66m2orOirj6Q7m
ZNRDX4ZsVxcZSQzt4K2C50nC7uc2ErNGOxw0Tf9TpG1zaewH8jSEVStNBYdJyazqcvk4SYHWcMai
1rtLL94GlhEMuocOYhLUrA/HTx/dSL7HSlIuzfmod0Nn+a6cS74e+WEFma43QGv+7k9ZB2pr0U1m
Ah/csI5Q4G4wwlWXoV6lIe3CycjoNS9wOWmDLyaiUNBdXNa8vUL9JSyuI+9HkeY7Gej6NCOZGo31
lWCUqCGJovv88w7nHA5wzOM+2DebQzwrsecEmN+5jRqcw4t+J8Dx+DPUuOYeTksttL/QhW6C6Yp6
0xwY253vdWQHXDpvSYDtReFbzGXE9SQ/G5odqUFzNABl532aY4eVKt9BgbSiS1LFy8rvLfwka4PF
sDoD5MCfDSZWJ2Q9oqZjMpJHAO98Q7QAvcYhyK2C2wWjEat+SMVKJuaqpu4vOa2Z7UkGWLhVHFzT
sdtRK/wcVsb275ASQfdgQeJHqHSNDMYqE2QdkCW2XmZgjBQkmvAkt4hFW6R416YqUvi+O0uFDx+a
09aXDK0+fIMO0x7urTORQ1f0wSzIdeKT/4vtcRQGOR5gnnL+Cr5yok493FuEeNq6ooo2UMuj77dm
KiL+ySFOCgYboilHJ3WP/cvC6xrtQyT/PemdFGfdDICKQ8al8HM5LVED7CytVFMEvj71xKpBUlLN
IFaIeAu0qggPmc6fdxsuO4kAuEE8pZL37x4VwTZuJX1tLXe6E3VFYHRekOJoCzHWYYPm49LIFQNK
p1xhwzYkDu5GRasYJFjV5v1rty4v6a8/POBhpaq9PEIKQ523+SUwAx08FQQPd1IHgeungped3D49
U0FUIIRmwia33Uu48mch1iP+C8RsVWroJVkhDeBeq7shgMS1NbPxx6cWYq2UPoY63pJonQBBSUV3
V71hBhFbVMnF6u5rZ9rExBhZHleBe5voq6LiU0BXrzDhYfwWBZvV32WX7cycIMswGWNNIXhXBfv6
QVavlmBrZr44mvEW0M7qEO57dtOoCvFPowHweMFN+BGXV2hC4xl79B1ko3aye9UaX7gNPk/YmstD
a28EoTjSpeCQ52+PWv9XVEIBIM+qRPiSNW73X+0u2zm4cgM50JHunM/GHF60halE6hL2CK2dIVub
AnTX65bsiJxJcLcYPAiiDxipHEdkHvC3ZmK0kpLp3aTvVAyzr/TvtgN5fTC5S/atT865/qtiU8q+
xz/fm5S7aDRI2M7FWIaWkw2KDALCcTNQjSzli+YFtHmiMEtidIzzuYrmaNcUSiNNcBO18VC3wtu3
q+SIKCLVJWpD90t3jqcD89XooC15IngzaqcdVHdgT7fEA1ssIKWZ5Ohw9mN6RabXPg7A/7qihl8I
83U1LSBX+BwmPCB7XCWLBVObyMswOwllPCQWezYU/naTJc9XzFn03yoo5lY2lzwrk7uzqHOhSEPV
AeGRBgV4qv/iDa+52DVJqqx/JDqsGn69fGGhZYrkVLy4G8DDM2c1u+EswN2Hk23VSUYdQT4usYjP
S/I/FKec0S35NpcX4oBxYaDSIRalsf1iVZcl0T5FKlvApqMrPKnp4atZwHc8P/eRZYly9TktO3Hb
fPdAa/8JS9O4mL0SpJcJOnils1aiyZfi4DGoS4kzOUpnDS+sqXtw1Ouk/+6IcI6lQyBMh0bj28YT
rJ9yUbq3UCCM0q6vkpjBZmOab8WbBm0RqhdS4xF9j6ZqDE5vKzCJm/+BPLRPqsN3UjKBrp4cPE2g
6euDYdL3ei6+tyuVoDIs+T3hSIOvBzW3mk6gZm1KF/rVHN/e+uBnrdW3pVfiq5srbHnfVUHoJxye
dqIJofX8bUOeftcEVOcZVHJleHM93Jpz/IUJoaITc5jPBnkdaPNHO8L8BayMUPPuFHZNJribbsjf
eACLo3ZCfqWC9hw8iUmTm5/OYqLK//Pgdz8F/PF4itCkyglfpnOsGzSp18xi9dUWMwkVMZ0phgrE
qk83gzHPs0eemjb1Na4C+U5+kFeWgz+bk0CpuoPhYYXyceyvz57IoDtSYfqRz7GEKGIqu/GAuPJb
D2/Y8EZi9LaTI+Lln//WZ8RGYJFMjlF7eQ+M4iDnu561Qnq2v4SKCdtPJVkt+jzxnSKppftkBXYf
Qg2OIrPsBz1btRv2k5rV46ojv02UHKHivoDneBle93D3UIC7tWcpqq/UmjqfkjT/Tr1jnheTacJe
NEHqaACYMwckL/Nl8z4qKKRG7qBMIlQK1Vf63LWmuV1xmzIl9DtflJcVWMdR97TqIcCjoPQhHtvq
Gl7uA2KDsxhC2NjreRpKzNcJnSG3LMFchKuGDbS8A38g//s4xS5ORCInvKz3rBT60imLeIH7jwuR
h01IN9X85UHnRNEAUQMMvjiI+xZ32KA7HGAjTKAEYz/YXj0/HlZLaamorJufCmVoMJBLAxkA94UH
tAVln7NIsnk/EpWYtX3ZlVYH3SAhvBqoTBOYa3SvGiuvXWSG9uju1RE804oT/FtJ9r5ORcW6wrt9
qwMQj72WV2K6upsY/RYe6NsFpmXGCGDCsZTq6FANmOHfQiwm8SUsHbkQBzGrdxE3FxyL+HhqbgqJ
T9EH+NUVIY5bEbrGcuGTJR7lBrZgwA7dFiZry18yUo+DQJXpNJZ3zUyTW1qvVlcEWUoz2jg4CdLk
jjIYqvi0QxmC1jW8+hE0ZhxWdkw6Imp+L3BZOzaYAoX5wYZKDYH/426puxEIdkfsACIUrvFeBibA
2PMc+fVK2dUy7v8r7WOSD7AEp4wtXOWGO775eooKpFt/71UY9M1TbNK9KlP36Ca27yTl6jMT/b01
ZF36o7aquFYbpeOnehawPs78b7WVLiVJW5Avg6uC9zfutZWJ1k8AJn3yI/4TdGQHChF+e+V6PMJR
QlBYll8944UZVScZ5L2SsgJOvv3YSDxBNx+29SrqgjZLvNYRc0RQ/PUzVG5Yxcg+EBBzO2MtB5OO
AQTsqPHvQwPmUpMxUjq5xYHhwO9NPw03GCLwjgSUEIig4G1rfDtPS/O7snSO3TKBMNvhlpQ8epj7
AH/ii8f7drkhlZbrKCQqzCFXIm5UWQhBWe8PuCwYCjyN+iUqqNEv9bw4GnmTUEvBLaWzQif5REPr
6QdIl/yaxNORF4UYJCKfp7nl7H93dMcv/ksKPnvcWRt7ZbC9a4OzilpJvCAfyeR1wZ4ecWatgWXj
nrJhrZIBEKKRkL6fBCiNQ/ZJXgO63ouSYEcoRp4agN7sM28ozyivleXQAsSvGSAQgsnI6LdNtq2+
pJ2nXj6Jrt8OmG3LxM/UITM+dylv/jnOlUB/R9LD7k8zV1VMwyf6o00QLveu5n8etqOavngyYoF/
N7YkQFIYIhySh11bL6OmB9lx8fr+m7YfmXfcZvwPTK+1ljPYerrqb3oou05oLxCVUnivRouW13Jw
qz1gG11RVmlEp01xWv8+v2TostOrLrAUku8Ljknj/DNlZjlBx2tZaROzfgU0ISqKS6xPN7KNgavQ
TT5CSAJ11uklEG6AchNpOUNjWmNZRSqqsNaSiQ5h9dPOOizTdVCQMlpRndaC26xCHusm2Gy2TeVP
VcTTwOnET92Zpl+7tKFUWqKfbLkeM5z/CTVnbMDzfL4OG8g0AjHSEJtcSkvLJp1fj60K5fIgWs/H
JDusuLJMduFnoCMhArg9H9I9Ma6V5vljZjYxb8PwaLIwDzN52eddtwLEtqUCm3RmBErBNLTXTF/+
AD9xaL5uezDf4Okm/Ttcn/wFE2KR754iBKO1vSRYNJreK9xGvaBaijoeGI/bsa6E1yOw2qIEGAA5
FfwaFw8Rj5g5gl73otSI3mzhvRGWUvbtDS6yW75Ld2OE74+/Tpcm8+0oMSkB40cU72Xy9aG1gEog
1Hkc3tZ/9ZHDro0OICM2JmhSmCq6BPpGJZ02J9W/nCpLU/B2AX9zSYj0M9t5JxS7OUPKieuELYNL
s1V/AE6LyW+NjlsPmf31mXEYvqK7KNA0R1KhRLTPP+iJWPzKNcsTcUYpLIwHC//Bu5msCyKOcGtq
WnzpVniIXGbxAfGQKZ+KVfgwZxx5OGYgzsFP0WUK9N70RJiVOdb13omt1McM9N/BT4AjbPbtojvF
svAh00yYCQEtnfcnNXWB59eguRu8KLJY1UpfHwT/npU7WzKzaIjdhevPre7fI/Tiauuc13F8kcpM
ewbNayIFylx7Wfm/wBtB5i0sYDZPP7n0+Xs+Lw3OWRdTEo29NrarixlWGDMS2R5TI8YM/5GV2O1N
IXWjoSBdNEWdqxaLU2PbTUyOgCi8g6mJZHeLRcGi+QsXFs/WUe1t7K8RZOm8LmQItpkNVZWnySQ+
5LtPbZOwGep1GtnD38ABjhdY2W+EaDo7W2Y6AxnDFilkEwP2knqfZeiGVm7/qTSQ4KWhXI0fxuHW
QTsa+3KYV+fzUgZW4sTcXYd50Ln/G5J85Fp7E7V3t1MVW9bB8f5nE4lmdMw69Um5Iqp3U2zvZ5xK
MvzNh9bcPSYrj9KFUN/jRx0R+77oRtwoTGyBOzZukB+tcnVvL9Vj+wW8o/9Eo3Ld7rfNL3VH9plk
91vLi8id7YLMu7SNsnd7/UOhym8KdpayyJxfc8BXQK+b2yljKSnuXeVvsvGP2fMCnc9qkDA2yXS7
+NGoEVl9V7+krQev/AuIMSifbLMWtaID/HgLIzTOq7nXE7rA+gp2CfE+sTt6HHeALk/QUDUayCZa
5pTHzRdYEYZawMldQUKqydJ1GTfWTDbCGR0eAJ8iSWhd49ilq3E8v5vvQkarSLLjG4vDSpRlXYgM
Uh5w5bgb8wKO+CQh9D+DM3yeEIa86ZC3j/MzvWtBOR6UJmGXy/X25TNdi4RoaMrQh3v12t3YOOib
iJ5ddedTi9F3l1WFicqjpalcFU/iO/meii2GDjT45VJ3bmj0sInXuTxJ+gq8uMZV1u4dvJmd2vsc
YvsXNIxgowQcJu5Hbmn+R7+jrzxfediI4BjJkFWaomtGEaBD28AmTwLWSe2q+b5uuECNAun8DHk1
hkmVRf9tqF2rvtxhSozZ7mg4xX4GY02dxYRjgcd+LRqY9+ulx9PONLoKkwQUrvO+HNC6pbShesmq
yqPub8KGO5nx65IHMjrXQwolQYIp/XVWrGEMDIALBRsIu/0bC9u0gMtKJFtCFjQozpaJH6p8/Wgz
Upxjl66bNPZxLAVs2R3lPLeVVtnitBNtEzcn+0ZRihvOWjQVUCnJssiE1WQRj8ULmi+YYSvV4NK7
uyxY+Bn9RM8tJ60mKLZASCcTrzDJANqWvAY0OSGRdgN1ElW+MlTWefnDnzevVX6i+6lzuTMK91Oa
k2f+6KJVwt+MHiE+7sYbofFDBk12BXNbifas24cHzOGQFLcp82PLBQ+pbXi1S2aN3UGQKga84O4U
OJlc4SrSw9PXhADGhfULgvNiYNDG/CwmdZxWBh0enFGh4tvge7/mKRPEOg82cuVLy3QaRuCU2HFC
GOJCTakPH1VZQN8gja54Rkee51lOkixGFEclWUW01Q4+Z8qrV7U8AwOO5Fv7KXlumETktYIK61rw
aC/JiOwXKdBR7BIFklqZdAX5lNOuOkxOL/KcRLTDyWMZR1dyJkN7w2ufM/0+qgsplcoKYrR1XDx5
I2eDMhjemaEDHE1yzxSCxuhRNumgB/AmCqsAt5d7T6CCvJDgH9+ceWgbTupP8b0RHHesen1zp4cj
ebX52MKkdq5wGIoQpAFEmO7inRQwz1tyYXg/HW4YmKNhfY4wTD/7d9xb9fZRUAyeU+wBMVI3Ddc5
Tay3rZDedJLwmejMZrwIPSma/NqUDiMOi4taj2pVY4HhKy93B4SLVRaW/eLKS32GgATSIiGuAPPg
CuoLpDviy833HPBBHpMf3hqpxIWIH48xs8hqkYbZdIHhxRlT4EndI9af+/rKsY9l40dXPIVNafbi
pAZV9AnSaJRIGSEAjykHP0ZwQ9s6We+ej0G0CVKg4BZM+ZP+8U8erj+9m8jEu6KXlmtBy1/FWLzN
nMx3ZkDArW2fsKMEGXoTkMoenAYkdt1akbgURB8NMXntmqq90zdHQZiqvtLBiBgDa+nUVzy7X+GB
gKztLIqpnaj2mQPnwFk62Gi43lYARGHsWgwDd0u6MA+FrI3ts1oFAqVcgY/ciho6EduNeKOE3R1P
6lj5LJegwaiNOHQyZQ/fubpxmzONz4HJUYoZxL5VsCSI7Z5br7FB9hHoUVqxbeugqqwG5RDG2Iur
96Mc9kw8+qAOf1jAPPHk9gWXqelyoX1HU6YC7GexGpsJ5dbB/8+cxEN9LvM+SXeCqECn002OlUlm
Ep3RDSVErv/qGikw2sSq+swj/ycb1J509kz248hhDJDxntLqIXnaA7SMkNz1lsfN2PDqe/EnHdpZ
zTWvgpytaB6PUy2vaoq3g/3CQa8RA6wV2f7ScIuDFYjv/ffD6D4V+tNf2WK400GoKxADJLhbfUbh
dZLcmDjA67WWhn18fjFhpYfcRhJgUVlwrhM1SXWRmifnz8yGMW/jErKwZq47s56PiZUg/SZKKn9b
B05oMUu+ArfDbzbQMNbStWv0yVAwNpve+hK/1CqjQgKeGNd7maIdyKqcYn9zL31d6ciIATrMkZVR
UEfv9qtNfKPohbIj1rAT874Q3HU2y+A1jU5hZYtClyyzyF5Wl9ib0gX0cxdtuv3lWDWATVeKfOGe
lORqSpM17jzPthFDlWl12a0ZNoEmHxh8OHMCeWDtQ4aA1vVsJNcrtTMZMe+LoErlafrnwGDaulJj
dOXTQYnIfAzj4iq2I2XTgMjSohzmJQbgR3gdoeyxCfnBYUoT+VOj+H69jxAcVrePTRk97KkKjT4g
daWAugl4K0jazgRVvtfa9uQ3lrRLSa5yxlKVuhCDzCG5Y28+GRXin7U62wb6jxgPfHD3nttFxGsI
YDCXyq0s+snLwGr4S7gS7vaBdZagSgSbSGMy1lCqIIDtDKUeE0Srcgcpxc1V9x9pmG9DEM1w6e9t
hf2uHrdVaVwibxsCN/5bDsdYyWUI5IjFxEb7pQoFlmwYeWb2I1oBhPhYsjOEqutq5gAgNk82VjUZ
zpt97KEuyRXUzA/aURZWd6lfrey0NPtqu99zALiUvi94MQDa++CAQZkDalkJ2GvaHCjNs7NTVIjg
dvAnIT3BF8dIdpGX5JBtF7LQh5Nf/cKgqonbrv0NiYX20SrMXzLVjXOmjUqPdOUOdDOp3BV8dJzs
HL6sK91T75RF06izOjNZUk9TDJADH5r8UHbqXsmATefbM7+e0EoyjtI8AT9Z+dnTrnZdTKUrYcB9
gW7UllcxPJ4c7YFHL/AUDXm5JuXpG3Ewugd36RX/ZG8EvEj5HHyAf6QFbOj3EEXvG9UNJlquVeKr
9ai7roa0iun6XUrVBd8+4KykltP0duKDJIGkh7KV7H2sYKO23BUnbNcPlBl17DeuRP+xByKI43A9
K4+xBbOxy+Vv+oU9wPznGYzeaI+roNITx9IfKxV84eN/UC5020DPxvrbNoxeK1scxwVQvP++tQ1W
WoHcrzI2FCl+PiWHc8eOq7fm4XDV7bxECFvhZrM64E3X20JJQSJNmkyyFj6Oqbovi+hHDuC5GVyz
krGPct51XfKGjDkF5yw3HD9YxI7z7TCD6en8h74WSiVwQXly1GbDUzUBxTX+E0Y3bl9VRvLjNc4K
QUhjaJDtyh1O3ERLUB+SkkYX6akrJIZJ1rnfTED0qo3Gv+uPPwcoHLPijcxW8HCiu8RxFoaiFbU0
ZMQ3BPCJlJK6/5Rhq09WjV3PhgOq5gEhSkzLe2gS7DoaymCOza1ngHPULgno36n4tqHGsWHiSnvd
uQedyyCiNc+Orsd8gVJLUgES6KFg5J20Utf9Rgq2iSe8/t0O6NFuSxOvBg8zNI/HhMopETEUzv5W
1IwaXh/O2//ADrZ5mRqn1BRZsHaMpmhUhapuNx87fhzmyGNEYJpaC1c6vvhWIc9MqnwZ7SOrwXD0
rh1v89MLRx0il2DJdCDf0QufGav7fetRz1GtlFwxn+yhI2XsISNt4Cmt8kW8dhDbLvEgt8g7w95+
9xe70pmEyBsgoWjMU2cQEhsvP3C3wCi02Dq45pPdYVpWEVS+GkNLJ3589WYro8yEVqlxwpfPsmIA
BeOazQIwPKode6R8a/iqDqefcX5cFckX3EqbhYfCWydq3v1tkxwERvYFFaL7GHWaHM83DrB68ph4
lCusGV7eE0TT1VIPawdmMV/JbeBitb3ZE974ccvRPvGuM/ty4cb9F21xueubYTSJlW7EMzyIzJoP
sEUMqM7aI8AH5Ba5Y841DIruKPs/1umSVLmY3bGydBcoWaV27cOr/N3mbkTlLEEA2tGXo0+QMKqs
odi+54qKFuOxqskkXKG0nh9Qzj+Miu1oV48xa3neJcTHfLzJuNwexGB2nQeI5ipZDfTX++aib04H
ZhZlSh2SHCfvc4QetSdeU8zKJgk+IjFvSOr7rwxuUt6hfFfIBcbXJYHTd1OiS/ymariWzgwFa1U+
xAUVkr5UjnUTDpox0sZ+iIxL72q0Q84KE55ZH09QLT7j5ONbGKj+zS5DqLdMh6B2dUKGQ0s9C8D0
lQ9XxJrTMJ4id/6DSH93fHJOR7gTaN4EDAcEEuUSfbxeji5Smn8/F1fLOguTvIxQvA25pk9+D24Q
BnZ2jh+P+sOn+Ah3s+oHyxaRgFF7d3+sN4l5y/X0mvvR0TCeas78jZb5EEfprbrqeZzt/ZRi5Ytl
wqbxcNvF+kG0wfaV0INngU9Wg2NIyAL+IpNHVSXNCkn8bBCeD9VyqjvyXJ6yn/+tEzje3/RGRVcq
GE1XYcjVKwlX6VFU0H/ejUOgXaDcSVp2LD2Ppsx5bdt+lG4qnEiVYPvEbAKYczw/gBLrMFmmtPuR
kbF8up4JbxuQYwbP1SRfYlSKQXk0n5MoI0PhM6/2XjspS47GUU4Osi9tZXK2gFbholQBvDtTxcYD
hFKI/91Ewvi4mmUJqpPNvedjRGOvJjeKwQsqFDKXn0iDXO9IHzXEXsO4FVAeViWZ0iT84WvNp24I
rppto0BHTdBhVfS5fa5ieFZKMH2nfqEU7/hzaAqmI7m4MDFLXeUkI8XMqbbm4b20Ehac9DJ86AfK
WnMHqs8T83vfr3vUeN2ePz4c7cu2khU8wnTmZo2q8phtTFk/A5l9hGvNl1gARE6wCNP/+FRJQ0ec
ObRf4XKiYOcMeNafIyEnQwfmEbVimdb28ReInjs53vISKE/sNvs6kXL3Xl1E+MuJNdzAJVBQ0MrI
mAv5+8y7mYUJImppj9jz9EV68UOre3quHogDu0zJW0H8malzrVh7L2ijZ2PGn39Ev09GaHeko+5f
+ODnef3VFlOmnN9GDW2WBLnt1PQbkBc6zG1xowA+kBnrTUNOM12SXZEJXsLOloVXNDuK2+HdCUxd
qFyHB/9KMqfRoJEaRB/tQepE3cQuwgbTvlmEeAW9lVo5npsbWX6MlR9iEgW2/ty4ITvaQlI3rQlY
OLk0tb7qTSJ72Ta23jbT9G876udrnW1GRGam7BLQ4/yyeRXDUr//heFxCdmj7QLAv+4lfEyUK4cv
9fcHJ1GsUCpVwO1G7qwmnWCaEz31btVgASWaah644y6x9GwiQFhayEYQQq80+30de35NlcAiHjA5
RBCFNQIkly10U4MV9SgJKQtU5kUkJ5cXs5PBvr2BLNSe8DtO00JKH44huvjAlrlVId5ffKobxFsQ
i1XrJdejVuihB8eoEJgYyH9ZPdKGjQrevb6hu9IS0qWMTlhLVXS/0zgDi+mbr6eF3ePJNCHA2kMM
f5wdYB2sYFXWdNZOEFywT7dL+NFDLUUxx90zxVMGN9F1Cvx7oHm8B8KURkrETI2AEcQI+OkQQ5HY
xOoK9btD2EROMqCMx3B4V6uCDZGNDwlLD/IBEIcz+qPyTWyDESyTuEOj/TwFC2q+Cixhbv7SqFAK
S/3ot5TJIcaPdtO1beSVwo9ckasrE9cGcCztsyEHQRL4FL41OJAaHQzxMLzprhHACiRuKgctkEWX
rgQ6rs/3N3Jhlw3s2fQEBnLPkTafG/dhnHDtKC3ARKRkG0SakcnNN0Hido5DLKUDOajsCsW4ejQp
L8jt97js/tqbs+qUjImbawzlb08psSHDk1yGcFo1AG0H8y9JLqwnKN3dTMzejYyqoISsRQI4ea8x
ScTUPRhN8nJRu7IGdIY3452fs5PiX/ffwIEexClof4U8+uAkQG3hDY6nzGN0Ual0K5GLao1UKqrm
XB3CqdDiprJMSaDW0iiIPIi7XkAGRKi+2+RDcJO9bAazyPW/y5fA66rov60NIDFURjLHzx/R+pgS
ZJ2VHE5ZK+O0zPkzkliun9QjQ0Fg7e5eNhDciouc36ljM6MFDtEJNWZKF6Qh0w4+S8uzU3ZCVGx8
lv8ujFxPH2nQU63kpmu4Hb+NfxPSBDmLYkncZ1nRvuEdjimc8nECbcj/W5ZJjz/LtCM2Rak+nIxI
lMFk4XCaJA3XhBMalyjlIM6qOKTtA/uXeK+NhWX5kLY0FXAtperQdHElzT46Wrqil9ddbAFVnsoE
c0PNSP3DJhdRljhLcmAAllibZSbAQEQ/aXwKm+2H9mfDRvY8+FVpf9CKuKBbc6zmSMyIWWpOLfnW
2yPQWN/B3BxDvo5TGMJvWWV+uh1GE3d5Fi/AYiNICV0jmdtLa7RlA+DNLTZ0DaCctRRKZXPU3eGg
lECr9Brg+23lY1zKX+naNQswdOvPBSBQEEYvwHnULmAV6LO+2qk36PqMiEheiKeD1/eEpesHbNYW
jidszmC/+lZ+2/8pFYfGc1R7Z8GtPNvr4gghf1q2V31GhbidR5fu6EgehNL+e25e6YQLJXgk40Pm
O4KAmou+QywrXNqRli5F8o8I7JxuAsI6OsLniffax9rY5uCjm7ney+TcoxkK9e0JSh7xjx2f7ZKN
Wmnwte1Nqz14ZdfCtM+yzHeKsJ8LRczO/YqlA1vCBBzP5bgrpt69JapeGMqgxhJZ9xJbgBHg6S4f
5KbZMOBibquZISaShUZYQAWWUbifx0J6uD+Q2ZWFQ/B9YuHv6F1/KCENdfbTG0MnF0b10QIiCUV3
k9qPz7TGEnpM8tAItoHJLgzsUjqneJm855PH3kop18JMteorTpLssWGfI6MsGNo/IyL0R5yzdjrA
oUmMkPHFMVwlSlxSFu5s+W37LqtwoQgZmgQXeDMYqN+XLYeOO59o9W6eZ8uGDYzy5r9wwgHHrJIC
eSQBItC3hwNGFI92XJjj2GU09PkIrqROLQv1fHSJbuMcQmhuFh+J3yvOn4los8VuHPkgVfO/Orhh
35Ka9yIh/KcbVa8Kg60+Vkt40X3eQ1U0GaynnBVg14Ygmwa+9RuEeLSoAZjr65IRROAI/KhzG0kP
a6xNjb20BRdIEYoXmuAcv+JUMAEJwHjKYT67151i6zXvQbxPvR57Nqu+hucO8Nl5rqbm7yEhB1jk
yWimij4fF3drGo8qddUeJTGl+HyX/8a8O6jurC2h3QWoAPOqAWisyTRi6tnkHaqziQnM4UGK5hcT
PcnPGcSeRUfGjZAnCg7ExURxhcSjSY75EA+ZkvGmFVajrIat9LjGiE3zgQllDZcGsP+USiGEbrpi
oh3XoetaLv7IeQm4LOdkeLeKf3YNjqVB+K5FsaDEXffObfDAZgGBaQwHjgfmNj5EvsH9SUZ8o0+D
II5f4WG/tCDppJHjVgfU7EYIeRqgvNGyLnS9EH55UjggFZ9V+czhqf6rwkNVzv3qtXUpi9TRsKln
vVtH+0/2CKv9Rm18aEacEtdSr7dM+Sae81W0BwlQw8BMZUk6S3UuIV4K8reKtuz17drG0h80Vhuj
pxBkR1z8dwaVWAtQfgKbayATmGT44UECXkQc4n95PKe5smYzf8OSFqfDa8u6xNC74Qky01uX3Er6
3oZEcJ2aZYiVwEWP7/xkp0pn3iHWKCNkazBXB30Ee34Y+8bPBOBelv3S4F6BVEtuyDo2Qk/qqApb
MfBYdn6t3gvHG70qrbHoQdZ93Qb9UhOftR7HKg5mvbYrj9MDltG426+/QwlmkosOBhryc2ypjtRp
0YFXUWjLfMDSZk7SjFrmflI0d5OvAgB/if+kPlM6dXppEFYg3f1D2DWWYuwGFbj2yuVndfWgf6Kc
Z49npR4YF7paPXg/us9DLH4lP2SNsmqgL7mkzcQCRO/treSrppu3/3AgqvionXOi0NsRxkUFQrvy
/Kr6f8UHQ8HASKOlkrJFW7ORgV8hN1vnBXFLWrOHvrNrG0QZnYN6klSQctN6aDHuntRxumg5GTmj
Ao1rfO6AIbroWK3ogwijF02pNdeuv5KJMw/tR4/syD+1i3ve1P73cfMt7HDdI6YTCHU+ksG+3rEO
IBxVerigDwQb5jcUW4FimVwpm27h8yPuLkX3FaelOjMBynN+NewbTZHDBCs6OIPCxK1OAyQQBNGQ
PDOibpaSx9KBXdOaqPdn9PDD0L10l4tAhBCV6IUHsChqAaqiWEana49mXugT/sYewsFi+7TNHX0Y
PzHXxDAbI42Xf3BI2RdPpRgDT6WtPs1C3BR1xulqKHCu/MB77xUoAtHzuNmQ03uLQ9ysYmWePJ2l
DwfjQtu1yCAWA3andGrHrjXYtXUi55qaeGBmRqES9HaPczI+ESsabyagMhdjmXGDrsyBRF3vGOma
CzJnflnPp//yKnMWX3d7z0sYrRr3nd9X+SY1eeYPHAtBhFR7LJh2drLNam5+V10vCs4Tk4Noc6Fk
GVFRT0U2Ab6nF7ORgRyjju9Ikvk+UAGRf4RHKrwlWLwGcqQYYGtdVIJ8V9bZie8i0A9qTccYim3w
9hD+qb1Yj6gTh193rJHoO/wuOHEnt3M1Fmp7qPhICon6HaZtHY/iJvMFYsBAZQ8qJHfkuWMy7f+R
N1bW5uZ5N+vjZ4n7WjeyK2wSf3K/8DeBs4bxOQ5q6vqi2Ec3eW1sHSr/GoLPosIh8igrhO2C11fT
yIOuGRGqh6zAAj9sYQZYjOHHUAUqjhyQV8ESVBx1aNVHpQBl9fn8cHDZYi4yFe5+7+MQEgtcm3r7
DA94varycVkBbnwCcoc/wrkPhHrnbTDUuaVRluS2bbnRmK7EkDYka0cNsYE+cqayIf3dT1ecb8+U
7ENo0py/JJPXgIxDK0nQaE8/pqEsZCbi55BvwaGwxdwk7KEtNPitwJ9+al0qN8KFK1CGL3aZn5GF
d6Xi+r357NKkhlHtPTYf3bWAd8iAqKeLrOuVYmfxoy9k4jffCHX5rEpchBpTVJUHAF5Gr3n1yaPE
9iSlCRqMVn3qE5dAxTR0JnxiyNjG6NXoaJIrFVXDoiflv9zfTyhyWYB6TWtyFPNIqOlFgnJOj3g/
baepD0G3Uey21Vuqh2HbaYGHJ6JUeMAjiDZN43AjyYZo8DUca+/3wBqcmjHu7ihd19iadYZgqEjT
fo3kaUWPDKOd0Jdq0+1buJFRGiw2AEk6ZgVzTgWSrNknE5ov61PG1E6b1iy5RBavJLbROIphJ538
6KrUBPUzlqLQjL8bMA4l4c5ZkuCjZHtFPZoK51grRwcv+9swaylO2pVCvjydRqDA2B2vQGFwHvNb
fdY7Gxzxrawt0IvISY8BwXYYqJPnRkurKU5hAZMANx6cxcxk3wevuqpT26kA55+E1xhsUqSWlse/
VxN9tpFsw2NxT5ABKfa2cfggNtFOvdVzAwuMSQ1SPtJvtNDwNUh5KZepPY0dsBsUNZM8Txl1YD42
L0MamRxw3g8DrN/1xe5enJ6A1g/BX+pll8tSH62IPBtkAILfbxvcFmD3bJkC7Tx8IU5hOhxSTxas
ulaWz9i0Yjt5a4U+mqa2+s3jlw4rRI4kFqTx4SNNsTmb90Jcpi2ZYIXfUuB1OhkQCi6YIsw518S7
MCveH2notkQr0Kg0Q38FNT/BfXVcivibY/kku8CDon/XAzDTD/VjRlN7TmjIM9pB+dn8fAj/c/t9
9WoObTxBksd3zm1jUZEVCLQzJlC8tXBpGsaBvI4QeX6czqWS6p6tpa3RWRNVkHg2oQqNnbEBqQxv
lsa5cJeO/GL9DDzc53S0PvNJXqaug6a3+MAQujkmYm1TBXMRq9QcJga9PYNDfOFA7zJdqHcQho3Y
3XcOflAEKwKuxVLY1ML+og80lLISYYCtia1IM+xFuX6KdTTzDeCFkPTHL8eZpkGqOB6j7fWLSwVm
KCa3Uv2ZUxq+aAHFn6mvaSc202ZB4jShAEHWsm6JRZPrUpJB656ONoXFSgnezQo/sfNAh25kLaW1
P/XuScI1jy64rxWK7mRpr5vh5oI/jlT841Dn5gSo1SSKwApvER9HBSAO4tsr2VSk5RdLbno4Myiu
jnBXPF7V91RC+aBoexgpyxmDT2GMeYQGaDSO/U9O7C7IlullKgm0g/hXBE9D1dyeGNEXPQXpZXWl
tX/V0it8OeCDEZOJ86VbpCd5q9I7jaW1726PLNLsLL1OZnE2h/Z2s+OBXrb3RzT9Gp8uSvoQIcJJ
eU8L8zlYRQk/AhgIfbbls35u4ays52/8bAbUm0uwMpVn+csIh94M4dSIQbzKb7BgZA0AJPA/LKfo
SvQ8i1goP8vwmr9PcUZ5NLLcJlkzyw+kzRv284Uh0xi8whhgtJiM2ZpB0NlJ0bXYC/Wdu3FbAQeZ
69JdvxST5le6hkSy8SBTWM74/elnOmtEH6U8RphKYX9oAzLzr2Oq5r7EmYno2B4NJuWt/dcOG+Wo
/kGXTujRXYG165VnvvJnRFhZbWqICbh9FI6128fNH4DybZUS4AGJVa1F3eQfbht99pkSbgiEBeVc
4TQSrIgnMysC2EoheuRT5UXxWCjAS2JOSXTo7FbAjSc4HGGDAYo5VPp1C69rLPTRNtkhlih5e7pI
Sb76vOQWmlIF46zxuYROhsj5UqHVPkHyNsEKkV6akeia2aZ+uZY37ZI4PDzH9MNRllm03UUheixf
sTKutJ0PzYVpfbSTy0ja6P+VgsJSm05VzAneZqzBmG64aFAhIUnC7awsa9Z2EKx5eMkKUezqEGfn
bZLQjal9k006ts4tAti7uDaX9ZzzTUQZMlzoBslPdIAzeNW+JLDv4yVccGuakXegkuVLrbIxe2le
8KM8NHNCFKQpUwBN7/ZND3Ht+ar+La1+H9oyRC6aVngC3ZsBYMfLwLyEafgnLGjCmjEHb+XDoBNs
4OAATXFGNojzBwXT1kuvrbs4Ui3hMRYd1V7yHABxWFUS7+5M6h7caKXfjfOAq8lm1OeZDK4VSXqI
86KJg8VF15j+/3OxrYv4+zF87LZDlSj+QKDqUOQDMz9+ZFsYZAaiCvIQr+4/67pX7M41hi2iB6pt
dSJUcAMQgPalVGfShxkosn86SVZR7iSGf3nBhGa49Pr42DELyaiRJSLofcwupb4MxC8f/OLDsDZy
nrbaram+LgwOdz5T69XB+gxhDfSqoyxfHrZQfh4lLXFIWOZX7Y6Iqj1Xoxo2RTmYVBXk8kOd+u04
EC2XDr3O05dp9QR8dXJRqcq9TULU/SIv2BZV85dLjdYUY0c3HijmMEo9t5FIJG0gP6PKWDlCVeO3
YY3nIp1qZbVRUHWQbIH/+mAUzehD40XqXWdY8NRidXscsJLUmzFiAMd73B7/9D1ZkeXMpE+vfJba
JMitX9fE3hwbGAQjdXNLG6oCQ1YQkFNw3l0d0p9aNgUGWEx9cd4/20RLGvRXwXTzr8OaqjmZU9Qs
mKT4usHmByLiFIxDH9h/fhr90MbF3CZxaXhvfLY1zddOvixw5UpVwMjr4asZXugN9ZuGxadeO/AS
cXsV7cOCbezrROq6zTB3CVN0gAAHHuLpySy/7fFPuQBbp/yUw+kGOWVfAPFYJbmQU+8QUkhqCg+5
rABFKbOTp7HW9RbeMo7vCgPh5UqVJyX62fivZYYX6mpRdxogLHPfEOzqYTx1ijr7QD7vKxueA3ii
2kkfHpobY/Gw6ByGRzKZMiix5XtWK+/UypWV3f7PcFCUrmrHigNQCgwqdxiwls4czJX06C5lS8yt
b7/o5LopIw51jd7FChGVM0ZmN5mBo4s4t41E2P7HuMJzSmBeYIDrCX4BDWXyMg8pqTYhZk05nO5w
vQ4LG3FRCbAAuy4L2sB7xY12FerCqzbWaf8i2RQo1aygKCRq7tIJTyX9GNYjrG5D/hZMWlhsiwyL
etclOxJV30XRszwVGYnDmFN4deSFKSzoVBlVijgeDmrgge0D3r0RJdQPXvM39keyKes46FSdR2Pr
WAEOyhz9dXGfIp+h3/psmPbK4elAlLeh9zA1LlripGUTRdnmuwBVdYJZQ5t9J6RLvOUhP2z1nenX
HJqJ5JL5Eqe/bHHHIByP7PKoVgCi+r7s3wjG88OsOaPqp8uat0rVsPo6qdbmPWsIie2FxB3iYokX
hf6jU9dtDle4XFcgHchBDnKk1mWyahktmXf1UwXcJX7WP2vEjJiS5Q7WSJQHthIx0Vt3/F/oZdfd
3lKQZRN31DmBY3tHAvEXoKriGPdXyrA1f1DjTEP2jaogtyMF105edju7uODOYuCm7/mmKq9bfF6S
a1LCq7BN4VwYCUSrnuOBg5/RpGXZDNkMxgZBubp8wBwsVq9SkYO+JWACapTrQ5sA7mOL9N5ngQUf
QDdcP7Jpg3x/jXLsBwZrrgH/yaxjZEvStUonQMJKgGYFoOe5Y1kwqIi2hBW9elJdsTcskXA8E/y1
jbr0ktYxkFkwabmXDBpQqxgMr0ULooVEDL6tExdV9MbWSYp2YuCQs2O+G6cHZQeXyQPnKXY1jNad
M6tnn18OXNv6ypT3Bg7+9MTo4LcQpbpTjitm9krCXDgYVlwGO9iukIQvfWrjCQehmpqPZ+LEQhTD
Y9Lg2LdpK6+tzUGnoRA2CqjzP3tc1rCIWEeCh/t1/EGzlT6rPf3TIkgodKQCGJpslYRc3xWXDcol
xwlX679gmkF7EOEFXpLtSs05V2Q+uglL+1s80YMtXMvczBKoAuPWaJBPHKX7CrapM5hYLJq1dc8f
WUYTVKJgAxM1FEUmzLW4LyZTFYeS+uS9GTq4KeBYjCWKARNEPxEZvjseIFOkhWbcqDY38DHDT0Cq
uy4vW8oEyE7j9m5juUGClJtoHeurRnLKfpfU6mu6qbsa5XycHtLU8AQYVvErjAu1dgJS/KJ3gTpt
D1BNbua2urZbEmuF2vhOocuL1FTON+lCnUCjC5dW364Ek/j7m344WsC6ELMqHfjIt/jMPiiWcGy/
MpkJMr1yomLwEHiZFf5WyLJYAGmdybB1FKLTPksEQp0mqGEGYtNc4/PvBdSF0tub2MvN6S8Y3c+N
E9SBuSj840i625A9tvUabWqSneWmOS6qTFmH/W/X1BEAmah1HPGL5U3tgo3jWti5lUUQqlY8pjdK
5W6r10XYjEB+5UxNdEpf6BYl2gFK2OO5FZEljxdNpc8L8Rm8kJqes4bk/kVtXDr3T3UDfIRVObMu
Qm8CnHDZbxe9+4QzhR8rpEFdftSkcBsZZV274mJgLQ6hFrHGby7LoA+uJaZTyUKcdcUhjeWJ4KDs
RfHgwfI7K9u8dGndz6DsrVsPDdnYG15ni1PVYuPPDt6rkNelU3f/w74QOcFS7B+rB043QBIAkX+N
nJgW3AEzP3/WZn8iOyzc7CqFUs0YESMlbtNV7ug6S4RwFeeMlnlfM10Oje+NQsvHTslE2b6MTmtW
7F+Ye43vAi9//csq3nXNikNKWJ1NLlYWIIW0NkhpaVOp2O2tswecKqPkOdR90q0VOGSnMZgSbg44
NENxDrWYZ9HHmi81oznF37C/+/f9hazmZyyO8gdFY4KpX+QzNIiDQv+4dWcTEAObPNUxDF2oZ7Av
Mp8Xy/SOQ5O36nGV07rRcVgKJdJ0sRs1VZ/QnjZkh+ty2BdFT58BUJzGvzv6hCXX7/68cO4ynouA
5wvkf+8PnA/lz8kpixAf2iy1LOGJayG5CXN3ian0eyxVnCHY+PUACdEVf0HCbx7k17WslRFGCaOi
HQnSMq3C3Jks4SdSJuGnRclkLm6d53mXX7K0IBxBb0NyOOuURf1QfbnAv6JmLQw20ReqJiZNTAGn
wtxJAlofkJ83C6/Z0WmdhRqdwACKGO21apeADGTmZBV1ZGZXswt+wpU6UlClHgKXWO8A2L343RKf
yAoGAhK3tpdy5FFjkgKcoSOso5W4Eg21VKWB/2HtNltvn5Gr3LeII8SYVeLVM5dUgA4siPP7BMqT
Otz0PkSAaMiy/YTWw3njpwNn2vMcM0JihHcJnaPInw0pgzl7CvvXb/RBwk5+IVMHZTET4n6mdbxd
RqEOKQExXVKd6r1zf4v48nRRRRK0y3W+KtPZnIYLbjQwd3RNRh4DHNM80a0DCkT98wnRbIGloS13
lAItLb70eka8Gc+dsBipgM+KhGIDgFgbH1L4MEAd/ZlUPs/bdG+6vH2glVNOJEEsYErL2MFdiw1S
/dJkvFJjagNK2xhiTMYBeq6KNtDdsxmSSw32e1fM/3o3ofpJCY71Hn4cFyHgBwI0rSrDA7xcrASo
3r7AnijWyfeuAUl67yx0q+/bGd7T5aZ/mqG3BbsjZIitD7aMDHx37iYekAJhWcS0gU6ULKVpEZzH
rldAywoLNO4uwI+68+odTC6biBNAhyRqy9BZcXSeewTBUX7n6vcnjUAuDgnUODY0YGJZ6ZjiXbNX
bwQ/bYHTikblpin4FIB/3Zvu2y/ny1bsof+iPU5ELW4hQ7v0jgM15lbqdzOgLZktmVuHqKApnbsA
GAx/8tLP+ichww+29sU1QN9wJvRtPE47ZhrWazmStAiKgwvYi/O31VgA+LavwU10DJWNLJ4KCWYy
K2NgOSMTzw07XddvredcF4miyoAvV0fSbLq1P7q4yzuC1LZ6vcVb2uMBAJhtsk542mchSU11o7m6
FBIPmaCib7fwXrjeO6oXEF41bVoy6lq5qao+EYzwBgssF+ySMzrMVCCjv7Ou5Bkj+wcXXTiZim4z
thfPrb+ylAwsZGEfmxK0MJVpN0WIOFsNZh/oSkM+bN4YI4afyAFRU2u7tPemHae2XgouXeiA70NP
Gzv2BjQiDC4qLOQ4lmFh1G25VFT3AaCnb9A1CKndFDq5W6ITrq3pEhNZci8xdXlnorxsUWRygoSF
LjOEeh44cupT37NFFXnQ6p09JolRpqVW1LwiEKs8/qHSfzDk9WTFxZ+heLIN3/3+Ko3Hmd8/1gQl
A1dp91pUHtON4qLuLwEMbxNEcu8hMhS0Zm0WTXZSUZJ/WrLRvF715vnvjaAYEp3Ll7+NrrAn8ysC
WypBNIEjuFxkELz2NHymi5h+o4LbWr3GCf2iGiHe+3i7DvY8h7OJDzqsLW69Qg5Z2lo2Omkcm06S
wcIxf0yqSsjgnQuenaTTkSvWhqmX7HnT1xnQnccRCs/unMgZJxXCLRTDp2KBvYLUHJ+GIDWWEZhL
3FNlnRKvqoWbdJUN90momIpr2q5ztRtNwKntAWWNHJI0b0tOlWvOiCe7srJ2QP+DZRxXaQcqcZIh
Cw3TiYSQgPphtgFstaEg9+UAZqY8i1t/Wp5Zh8ucM9g/QQ1vm6B0oakZJLnbOccILhYvhlvd9Acm
yRNB5etmyzoWuJcZNRv7vFimdGczqVXrsXfWq2J0TfPWCu9cXEBxKj03OZzIdCABDUYh51QIhHqE
L91QDsPROT8V5g140dJIBBtugvcj9naHpWaerxKrh2mOsBQ8/Ceg8VkQFnLm5ccTqiaYR5nBvu6n
ayK/Cwmdcafd7BkIdLEtArj+e6UsPhATyOhiwnn6Up074sfWvoiU/HBJ3eDq0qHIxuNawnjTD4Jq
9JTyibDxlYw7semaP42v4NrmK54kB7BcvMcPpvlycBrNfa98hHmrYgokHn9wuXlM8XEalmYXYX+N
er998QveNGPLAqaVk7qxyz8C7ACk3PI62wW32gQbvtCPSIMDcUNMZq1/DTiT+1uqbPJjxO+xpEzD
IrO7k+WFf7KTDyGwcLm8FmiR1bu+lnnmu3t0v51fOnNU2gVd7lCfy8tVlA8TNpVPVKUZuIdFNW65
pJ2fC0KNPBH9ktAuwI9AsiAB6w464ZVrAbr0lHA4WfY4r9d51E7WdBlJ7Zu2JJp0xDfKbyGCU+43
Rbt6LGd3ChV9ZUyba1LF+cpiFxecnZQTeJw4eUA9ovzABiudoS//Kfu/PwbT7zkbb0EVL5KRDhSF
LRgt7KU6Ee/U6dzGLvN3hjILj+IliSu+aTzweAXrKyj+ZcKP/LfVpPyCMUUlwZ2tAeNttjG6PmsJ
3ZNo8mUDd1kUkipg7G3HCXEcl0MsaQyeOBCzJL80nT1MeBYARsMvffwSNZXLFFRS7Rl8O49TjBdp
0HQ5rwd3ViybnoAcTTJKINK6CVgJvkhUmMiQLzKslCPc/9tCS7nmP8GmtmXUzFK7+UYLJ0erlYKJ
jCNZkjKmeC6AmKD0KBXXRoSJS/swWfTxsKmLrzkuAwNnHnTXTib6vlACH/Y4YR/0Nd56qjlQL+M6
IQuZISgqIpMZC3WKB2Xrtr0K5OYpArElF4h2cvZ9P8/w/HagYCQWPGsKw+ZAZ4BKpZ2XJOMFTuaH
1a/nVF508Fg0/Q+3RXoLYOlmeheNqBnUnHkgd2iLgcrMMycU9p4/6R8rcihKkG0jIBrFQ3qsz4TC
dUHdJxgG7eUvbRyFWTGbJtUDtyVRN/YbZ2gxplZjLZm9u0r4E3QjYNUWZ02dByrBs960+Ul+YI8U
sT1Uy5qmhfizQHOS4WuYR23Fw3d50M171s0foGN1ToKQUJNvqRRyOw4SWxNK2ODYond4HhaGb3do
JQf+l3PJeh2/jcfXOsVXTlgWAkIbOZnUomZN343h7emxH2EnkktSCPac7AcNRYCUBbuVJmKERAL9
Wk9ndkO0B4KcfyKHwazouk8UKqYhQyj6YwHp5oMaLoY9aWTz0CH9Ukzcd8d8tz4s2twZgLRyXOQe
SWjahEJqX2dVEu7tUaGanKPXs/asNlI7cJyYzT3t/ND8yJRejVMJGb4xL4ng0bNP6ET06drGmsDV
ZlB2jqHtzNKiyoQzbrVfuVPxExNbKif2UM5lIge3vbqZyDguKF29a5i/rsu7aoK94vIRZLkpgIHw
riHCwoRkFUu6cq1oKKWDoeLg6YCuYNDxfWDU+IbOJAfX/0HhB2scAROxkGm5iP3zJPmQKs5OqgPJ
2PP0h/BdOGTC0HIaG8zstKA7waawnI2AkevKUAb/3LpHPOHIr3xAvUG7Kh+KRA+G2XCgw6lXKsJ0
JFh5SpPqfhfKRI8bTlsPg5MlzN87Tz6KGKK/o2zSQnGummidNv85nn6KNOvhR8QlTCFHAQkn8hc6
qfz667XJjsMHr9DCcVq/z2zYujEP6CCj7kH4/ky94olt1xUs4f7863G4yZVk6R1pgksLhCO9gNKS
3TtiKwMnMHE0a1YtgwSwmSmhI3YbKPXChCHOYZMwT+y854kzcgxT6eie48qphgdl35wm46I9Z2up
QFbtaD6qIG4KPq6GmUsXdXL0aum3IOHWo98atTjCqhMSnJdoXVp+ybZNCe2n+5AWSJlevIqdX2GJ
a4ElI+tNWiNn2B86q3ngRhIrx6UdIUXNz7VwEVxrtjh81zoLR8DasSlRJE1zPHorRcyU4gaJB08q
xmkRf46EbjGnf4iz6A5mR+lb/Ryw0LcRXhSodK3Ys3oQ2dfSraKqeT1w2T5V7VKGQ7B46KKoTiOf
RLfNeOOYPGjDugi3YgbIDHZ9F9+AWVMOLjIW5iDxRsukRmQma4F4Ko1gE5SO3qd5K9blerg97thB
c+Ej6iDvQvzSqEqTbTIPQiIUcrhG+D5gi0die5L+Oa0GSjWQyD87D1pf3iMhXmMl+sMCOBTuSrQO
OuRQ2Hya44MhuYkwVkFc6rbB/6EskdSfzqVD43KkcVOanYD9RRTUGrXaBLImRmGnJS8BpYHM3PLm
x04lVU4HqHpd1n9W2MhbQqSNInNUlpqv0FFlVR07NI7mXlYeMpSTlygGvEMqDHuq6TBSFEcpz85P
USDnC5PfbaBHgVj+hAXa3J6/UvTQvvM6ppfYUHA3Z48I+jAbQiGy8kbXLmz71uE62HuupuH2qRjX
xq3A5mV/c9r6JQWg3qh4r3GzrijX0WJtX55jyMQSRb1YjZz83Eq8la98vGWelxSfOx3e1tTKbtiS
N/QXyp6uPktqUYP4mXxuBd9+iHXVdPt5sA08evW10oJXvxb40+sd24jciudqwOuplWRaGmquYujw
rZ9XqrHPPu94ZDbZTmCcuvyOmSE4dtrLIEixJcsBJilx6buNtuwE2BE2ohzxcyx840Z17oK9f7OS
qxYmEy/B35IDf0MnET28ju1LXLAp8R/PO4ycPWtTuTbZmPniXli8M7XVrOHEDJRnqvvhnB+IlM3N
AzLceLFvr+EsoTRr1zziybxxDCYjZ+op6YlHRLIyt/1KgFKmtpaWrtQpGoHiSJ8u1L7EsV6HT9X0
H0ujwt3XuXOf2Bd4brrc/lWRWh/zqtFwEdUcqdQllJnruja2FRYMfMR6HFcygds4gkELv7XEnX7w
4Ma2Gr+5p0u04QER6tz2l8aKCdp4mTkBOuNWFvcemAluxf8gF1Q7CF5s8U/i475ibTBf2V/wSRQ1
CygLG8dSLAL+1S30BSU3Gg1gycSZVIhlohBdSEhRlUGuUE0vvji8dHHS9N6BTOL5w504jHVg+bvY
MHkv4ZCjRkcvJKtDYKqzEOjeZFhzGywyu9Tcy+mhrSiAJKw2N13wY6Z9J3HKN3iUzCvXgtDdOWyp
z/MaHSLgGAF7sRJMHEa6VyPLZFQSVfv4CMFtz6pI5/mC+SuN8lZksPEjfEMXQnHngXbG+9z2wIJk
M3oN6cN0u/JPAVSE5QBUbUm+1oIrPpqHDXwlUo+FMB7lXdgFluuyzqf2lgE/sQto7VQPGsrHX3AE
rguF46AQYGW26nO28DMirLw21GLeTTxCtRCBYRaD9WAgodYO+aj4vVK8OjdNGhPAYser4R4Jvp6f
UZbU14oqvxfW7JT9vcYU4uMq1sbJRCCIWBeMo6zOO6rfM39J+5JBKvXnaS4lCic2aFrwdVcY2dY8
aT0PiJ/h0oZjiWdcdqXYf/81/F8CBgoZzLJuzucyrfpoLbzzBZAweTxSiTAvip2ij7lxia62Nozy
vKjisI0biI1C5ffzhvSXDV02sybrDPIRWvYZ0rIMKiWfkZk3TYUOnk5KBc5IAhzssoysNzqw/yaQ
El3T9deuoG+Bs6yD+WsRpdgWcrqFmkyIK7xK/AMVa2bLHJj9PbOshSJnNX5QZ+zJBHlTpQ+LUQqK
Sge/fBs+2zGjOMqwHJsQv9y4AyO8JhaE5JBS4Ut1Bv6K7K02G7W+Q9u92255lnOA5gzt2mkmhHKB
Fqp8ICo0oF0qF7Y63nO7UGoXmOM21czaw3tkqZ+UlQEc7Fbs90QfSfcMYZLpAbaF2fvpVgxjcSk1
vqBPhzrZcXmPjKeHdEwJljsIq8Hx9k2t9hrqgAZxo2ZIbaTErvqs/4Ip+zLzZlYC9/wmdU/mncB2
hflogZGFYRH20WEhP5c9KJ7g+KBMOx3lXJugjzND1HmZKz/D30xt/NLYzIu7BSE7MqW8554dbp/Z
TAR834KNmS+6YezTsOh1mytH7YYXvtKkS841TPBytchCVLcaU6y1Ekjhhregasr4UZHJ2+T76/qe
2U3wjdsjBR+JIB9uVTGEWVsIxPr/KrR8B91WG+RyzOKEmOmKEABq/i8+MdvvpW40LqubENWWa81C
LXjTPE4nGFvbM5pFB4iV56H7Rrz7+EYM5b8PV5FAFiGQmpz4qjkmLqs1CJ18fmkyJqbirX7wPQkA
QgSyKMdZy8eONDz612XGc5eObw7uVbAYa/NF2ka+rqHwamCjyodDw68w7TJAqdim0wYsiNgUadZ/
FSC/zC1FIeLJms6H+P5u7S8oEpxde4/pn3ng6saLK927V/AZ2m6uQwOmGjQxwEABYFSMM7hJPOp6
xstA659vB92UVYodx5IZwk2Jmbi8FNZon8ZLDicJ5prGxSKPrJjboVX+GcxCh6yZMk2nC5qT63NH
w1x1fC0BQV9OavHG0CnpDizxJ9RSvRdVf0iabwPG46lj7MU0eGRxhpXmZEvcgTvo9eu7Ih+0zQx+
24pik7i9ht/SZMPb5e5ZfMrV3VZUtXwjwJ6p7dCVfEMVwpv1AaYEZXf3G7uPGfaAkM7Bxl8Lwmuz
6pTSt2eTQ/SevEPCplEzmmUr4ljk5L6Awc1iGf8NTQRAnjOk75lsEWR2pirx26RFEJJ3Z7q8lZVs
OxNEt9PUfYvZ71muAN8HREqTjrxo1P7cgek6tkAvDMoo9mtXxLqCVi2UznfP0cohujiCxo/eUgnN
/mrOt7q61ZdbcIE3Svc7X/1n9c5GmgBeyfVkKiObT0cssELT3zMijereqIN5iRup3o9V4ZAmCU6R
sPz44ntU/IqW9WKgQ1mCGCk3MdIjMUZNpwA2KLev9VhBD0B/+UXI72U9BakSz+1C6A+5IE5V2k9K
S/tAhRPIbHaK5KtuvdUkNJkc6EnXx5APA0BK8AWa33+OskIHK3Et8cgci3FiisUfF+4IabFOTn2g
CJE0W35wsA0mQ6IDjzL7hsPXd9EvNhD1ymn4MEmr5elvezI6pVLDzuRCCSOauzdWq5nPQe3kHGcu
9m1+cMT4peoqqjTd6SAgzV5MAaZ2c/bHiYUQLYEP7/lf6h7dyFfQ32di4EJL5Ib+ig9MuuZUtt67
2q0s+DxBswHya9KYlYR6GGlnLugeXVyGuNuT1veEmmoYUHzAOcJrPSOe/3rS0+CRXpd3RK9qn1wP
SC9ta+Yq06qPLv8AdB4aLOHJ+qOtAGLgKjLDtRG5HyEJzHsuFVqpP76UaYexS7nV72vyp/5Xl/oQ
6RsrTop32vFf3R/7GwIV7WnKK8Hxix32s9pqFbRCMKuBnjd5gNEsTkqe2FQBKEp8j/JvQEM0F8qi
dxQGggYxlTfi2S7wEJywuj/w4VheMjaVH/n0gemaSdGyaPKI9qFpU7JhfN3lPk7nfhqACfO/RnVd
2RNe6x69hwCmrs/CvJ3pAfFxxRBDruTSSpz4fuikzV2A76XMpsxR71NlYM5UCafmNUjZWKF9lN4/
104t1DWH1gvFFW8qiPC9dQ7FCGW3W6CPXhrBUUh9GJXV3ooYsOfl/9dChtdG/VuKvRGX7iMjaRGR
/GfdUPJHv7YZt2M39GkpazN8NV18AwQ5r6f6LhpazgL3UYGznoBwk4KXGZ2BJmsLl7nDpPjYbpQF
8fEY4lfRl45mWtfGZxvHrQ1yhlkiQfd6pWGX5H/HdO1V8MYVYfEWnTF4Q9tgv4RJ3FUIWFucQKNa
5qBuJCwl+p/HLZ5nMVMYT8orUr5tpqiqfvr/DTj/dW7VqfMPyrWgitO2j3wsbPDSgVWEhINv/WNI
059pf1//UgMN6kfJyuYh4+Nnmf2uah5y1xJlPT38tZODCWeEEgtMF2r4mH4pW3RR2QGAndJjXb7Q
amAXjZYgL4KYVTRrxYhZTqSD3pgbjDwAVVt6zr3uCmysWxaKQdCHYHr0st9299MPbdI7D19frGMB
JHcWiadrD6Q2xUhQ+KdMIhF2+Sd3imxh9pyPPdzG4Ao6BqK3CDih8sQQUacoyjmTIbZ6h5bhgGdD
8xQYPkXDSfQPvrIyL/jMmJXazInjmPjwz0nQTED2Agm7fmX4d2yJB30eCKAhbu4qY5ifrZdiwZWj
cPRz6b8mjUlIEQT1QzmOEz5rdH2PaW5uNS4Nxc8O0+FRUv2a8k/MdXjVBG76cwpjGCWqm7RYyHhY
asRyFbAohmrJRKWTGfnZDYCT+SKaCPv1A5d5MajgZ9zSN/APEvtQo4vmsrsuLKo/dDtIVCbDhvKv
ragcMUf+Mj2j5WYeqskUQgV3J3rNVGNtrICYNJaYKRbkI5t/W7eyeDhnR+5GcjHqBhG27SGxxjaU
g/MAJ9uUebpSMck2vix1p759OSOSkC+7eUq4YpAWgFnFDDfTm33iPn6aDPQ0c4Pb3RxpYYVF/aBE
T87fpXS6zIGN8puV2l72E9g+Awqb3CCeQhMgS4CXmMk3/DTqabGwBFVLuUH9oot4sHlXaRi4L2aB
jUc0ZPRWNBlN/1mliJZlLR+CrgylLaJ0HYgYDgOfH3hifWkn8M1c1MZcbFaIuVSGgpOZSAS5toUe
/+Sej+aR3h31douZjcsbN7U+FPkMEapnyXjW4BrkzEXjkjylV4rLJTCvoNPHTdsaCuUQGOFZc4f1
89/HyYRXmDkr06/3jv9ePgzx9Vry548peX54tuEM+NNR6duk48Qe5t3192MoKJQidxxj67aLOgw1
gOLH/JJa0KwiQYSwPMcggcyN0E+vLrK4ecw99Oacn5LmR2T4dW96fXl9Y+9XkQ6ntJDjxdOyyDT8
eZZAlQhxHt0z05ZUYg2sssGxU3hkdsriNjy3Lw5u9u32n9OYpRrtQK0C5SVbKrKNthx9KKh+oQbL
uIXrp1zPN7Wucz6aakXIXD+dGt9zzhT+WIR6DVLkIWzKE7KcbSmsbdN0JMZXbVUC0xjXgzlP+vRp
e2lLbFsjG4mt2pn1yPXB7U3EkA33lsXNlVW8R8D1WlGMwaPQPvAKV2vL1ITho85+crG+apm+miw7
+T4/dLyDTfUMod4NDGZWoEwpzCqJjCcQrK1sQ3oESNWyl+yq5AyT273H7NzFBCbOHikeK2EKTUNS
fF1ULZFCq08BBOKgYiAZGwJlt1e7HRxsFRbeScSadHtP/jWAbrtSsnIUWKGi8pMCtc0o5ID7KFBU
RTEUUU1IhHZWhfQfzCFTxppXVeD0cyhEin/VWtgT38QkWm1urLeqA1+SW+dN6Cu1Ct078QMp2TLW
CZ+Gbx2Fl4CUoI+qpsFwvZnKwc/YoS6XWAlGKIH03QrO04yu5OhPsdu4KCaA6UPJWqeuoukHapJl
VnoOYoDZ+jab8unV0Af+abY/FVONMf92086CCrJ8Wvh9YdmTDh160Hkhz513842R1m5aKoiZQ/3S
M2jlvM76lhnZ3lGH2QeKdd+f7MI8x0V7t5EqeOSuJIzvx5bnR2A3NjHB9UxBMHq+AC2WFv4DYXKk
5mEy9l6cflYV0aWAFLZpxCaI4lqjCebREseNBjb68pkfdNvwTt7i5FDarpRI6J5It3YuOpK3Kp9I
eoOyyUn4wdd3t5xqgyYMqO8+sl6iJ/JOEHwHAIldJ6rQfcCweQRWDx5uabVFacX67b5DkejtMCXz
z44UQ6xE/4RL8VfE8OJDHWpb3caKz66dddJMz2yYWyk46sdgpR0qeDb1v/ncRdSsE6hbB7scxSpo
zZtEGLiHzrwIejgStxgO9XCpGIjurCJJcVPnCFkOa4oBX0Uh/IZ6wmXg5mwIklhT/eHnCckxRG9Z
yZD39zQftBvOwIQOwKznt9VitTCLynkGvMKunkM2S/j6Yed41P803LPZ8JTuzt1UFqahfYMYilIi
EAd/vYhoMLHIvDFjCrflPq1P66iazgCjM4MwTozeCCAZ/pW9evyy1050n3S4nZZc0jvMzPC/RoHK
6r2AU4Ek5IcWcTOU/FIaEhtVhfel+lyAGA52hs7GSoWzzKSXemHsntYj3jjNUMUyQu25fi7DHVzl
bZOuhpKFADeStvjWMomXJD1OKFlxm0v4k/Pezj1hQZhnCdOJDE48Z5+2k9fIXP1eBCSADyIi04vQ
PPiUBd8ZwPTeeWkrP3Zd8BOPG6orMbLuNLRjM7HsMCCT5sjIMiNGzt+lv8OIlk0SuMCMr82FmwDp
L64ByENTVplPJ6KfzwL9k8UxBtl5pvLBpsA5C18TIlo0vlUXbUGzSD2Lw5Npwk/6ZhqFTmB+n+2/
fzMU3wW+K0Q7tA3WRM0XEJM+imatIEG2VquJdUiv01HUz8UEXyozK+TDZh8iBpIrZ+nkVh1n5rOR
3oAUPVkRgRLOtaYGBA/B6YXR1mx/9nY3rjZAR6177MmznkmRQQeNOaX7pBLeISABhhIhJauC5vu6
WX+GADJSbUTHO9bieOvWqNkTS4qkZtSpeNCSIx/fBqeKmNdmxM23mVJMp0M0aGqLpH36VbMM/0Ux
fVyXymD9aWxZJ6yUIY/0GbrF72LbTQ5/VpGzoq4rMwA5GDYzhTOKJ0XqEtKc3r5OBFseb7PGxYMn
cBKp5iwblrvl2BrZpczynryaCSyTu2DxibRUz6YyuH4hzzIUMWlBO73SRLXxSOacmOo2RR6UPmKC
xcKIRV4vC3cjeeg8uKUhq6z8RGl49xJDamEHEhA6/k2+oTVtdXcLq4RRLQJUUSPzgNK/CeoTvLk8
bvTgk+paQ7CFo93aa4MODjini2jCUoaoW7pLma+d62xB68D/JBB5hk500VacU+nBWzMqydB1TCHe
y52o28c5RWMWdtkHiJ0wwfDtFSPQTu6jxJuqeiO2OOuocmK2u9n7YiEat833KMsIl7UUuUrVyXSb
XC6M0dl0Cr5Zg48AwwKyoAuccQ7v7I7/hQrpspKbpDZ+NMGWw6J+1p/mioE9dAXCQBVy5186ajIU
/UV5D1xfuKe9bw+i7rKXcKNNxjrFs/vrEbWvngKo3BsTs9kQrRa4jS82FQzt0SgHRzQrKBzR+6k/
zVnJf9KYYXVqzlc1jNa98oAK5DIQ9Cr9rEcfWVoBdB0gZGtbj6Ho7JWFcM9rcfNQhnhP2MYHxlo9
1o7WcL4v4cD4snJa9SiRSZk55ixS0vymVFKb4SA9E4vdceG/eIgKoia6gDCTg1PJtdqTCtRHjDsM
pydb4ZPet4vHy3aXsFpYppziqe2UBaEOujVqNAnoOL+n22LY4XRM34CfuVn7RznGWbe9DoqYt57o
//1tlfjlGa6d8SnPu0JoBy9Z5e09EdSGPMefpZbfM0UJVC0DE10ZZ6FE7koPq+2dGQEJGPq4BzpX
J3R9si8H9SRPVPztOyyTCC2ICtQGC1RFvsfr9hv1x/fIQuDaGFua8j5Eth2/z/8YszEuR4rTEkS1
OQWb+uA6vF5prI//r9Uojvc/PEWypFYw0fyYX3AOQ4axaSlozozRWEzmotR4pmtwd0lBQ6LeYXXD
CZXWo6AM8OXHxkYqEKqs/TErbpMNB6mQoDoLsb4elr9wItulTrWh4kb6OrP3EZVA/lpUBbs5Rs1W
xbsn0JQjzDlBrIEIBuAHQUkuT4k1ravwRUYH9BQM2C6wOC/2AEBOE8XFTYvGoplqnDQpzBTtdhyY
XhfnCaqP2v9PEUAXwBhXUurXX676dEBc7FPPXvLdnBjLHplYG2ZxmMcEiFCkVyDtUy4OHKTC3MB0
JbGkm0zFmNAREIrSrCBIJ4wDnZWx7eo+uybMD+ZBJsPpnk8neTyBVio9zX3vpAtFFEtSZs1iRiqk
9+Hb2LVtEEgoZQ9woLLzCSchfnKyKgv8cCp40n5u++yapNJt7hYU3uZLQ3GEGLi2p+FnHGTkJi8r
uN85y02vv+ZI4gtgjAIWH1EXG6GhVC2FjJ1pnrriUx0EcFj8Zp9sVc7PxEjlQ43/8jd1GXdNlhB8
Fa6iFFLDcmuTlE05jqm7ZPZ1ovX2hX733gPecrSJRbg1nf71o6kHjyFhFZ3kuEzCbpNazO+SDBWS
40afoId4/ImG2/L29FybU9BrnEHYZ1/qHwFPGJmujBepIWYLrKLcoz2PtuTG8SzQSh/S7QfR83u5
ublTWqWyikXA2qeoaNvJgQRPHBxexynqTAldIyR4wCpGQuX7s5QAFeHilgDBGkholYJb0vOv+u88
KqP2780mbPJ0i8wEIhb7Hqh88/zvIqL7Cl6BCYAVHiuIu6FkJZWFPA77HjhVvwluI8ig0N+pVuqS
ZphoZLCjWFrg/RSwK1oIfONzY0yK97InjEHC23SoOkHnn6vwh4q1hQjKWhcyaM6fSdsQT7QeXcjE
axRSlzOniS6U1K40lf1/SVZM6pXkz9AMrEY3R5v9gJnFxwUZl9T19qo5+MuheyUQ105X69g0mhUA
DTwxzpMJTNZU8BQUtTtiMs6UMKCbFPjETC7ONWVg4WFev3r3O7QQVbLpXi+0Jmu96L4oOqZVxUss
7Eb9J7PrzN3k+oAsjMOwsPd6lq8Qb9WXnxmfTxYPH6qYkx7KY1j2q68YWr7vYiPgXvIeX3Fo1M/F
40rUvRhTdfNwkSrRCiy2ipJALssKyR44GWBh1h1cRjWKvfwlLdzJqdG1eN+U84qKKoDoV5C9QJYc
H1iT36ug5V7r1AANEkG028fyhgqVjCtSi50Fcy0Ls2SDInCNtmoAXnRhGYob3XaESebjDusCPcjh
NyMqfIudmNGRVjYIBSxdgtSPVFL4dn0U4aLmtW2QWLxxgj4qynV1IM4s5hIyeuxmCEu5cTYjmaki
UA7EFTsivJUeYfNP9M0e+g+4Kp3zgtEH3R9p+crjCB+u5+/M8CV3EjnvOI2Z0Y1dwAK0Y+kTL05/
JRKu3uAWeVXVVT1TLREDoSipFDOr3cnJkClvfHoZk7m7AHMMVLzaswPORiXMwzb2lDt539vbPPkm
5nsSW0GtBYiE2h3so0JbdMwCaz4kQFLGBwbTLGfVwtGa4n/bPLfxYV6ctDbrQsXThN6w2Q/g1l2k
G565QNc0pU64q1xVlWHQOgl1bbOS1Vo2mpnngO0LmUE6iy5AfPyXYj0L6uVLYeGw+uBBbSo6s70y
5Z09+SlTxaz44Gdd74hgqFAKWbDGc959UlV1oGDy4GSyor5X9zZtWMJVwtRtde7eGk+GPsw69RIg
zgK0jB5v3nZ9XNiv/vdnPvsj6BGN6onlFDawn232Qv+SM8kzkdOnp/Rveo0YqeALcq5HUSiaufwQ
15sHvB9SisZ5mdZv1Kh5SmOoRwI7NBymunTLbgzHRh+sGhPKyl8IjU0r6ov0rBEcANRWX7P3ZxGu
XEqtu7I0V7ej/3kExthsgxEJwxPQcjn9D8L2omz6Ach0d7+/2Zp4y/iTD5ugfrAWqQsi5qcP3/XW
AAXVE/V2BE/OwfKUMqsqhJeVO2+ILE9q+xWiKkM2tWa/058drQ14RXbXn1UfYwDrIBtZeQtyAqPn
9ozIZaR0sKWDR65hEfpIt85ecs1Tbkf6fv6hypKyKmk9jvepgeSZ2+deS1S4cZF2n4EXAF8LLvRO
HsC3xMAt4fSh/CzbxDKWunMwc61N913AraLp0U4SB9XKJrOE/me46TVXhC+SDwh1v9ceayKI5UoK
XmmLMeDuZ3joVDsn872ikq3gMUI0O4X5wjLQ/C+wH7TXgPQtcSI8W3j+hB0C1gv7MKv+k1Fa50sC
xsYUy9E6qCiKZaqIeAfc4kAdjrgrx9ptkExOSajuls/0+AGneWO8/9ki21QouEBIX6zkHZXxU13L
gcWR/UTbJOk8kG5CnGp9LtsAU4FLlGL2Ke922JVJXBOFJGV988ieNpKe8DiTOSgcHkP1YMqOfYLA
LuxhHDLCTLLvz2pxGPGmTeMiu9aPsNfK0B41dVhd/7wmrBd9W3J97bdiqO6Bd2sCnooDoIKuj3Gc
abJjjb+/70K1Ck9+2FVPphLY1aBklUlSXs/qCJAHR4qfeCUJixVlbs7F2dNjoq09BV9m2Xs7HCIj
DgHU7mrz0yCULjHm76nr2z4Dyzj9tf/ZqSwtRUXgLFFP0VA8W51UZYEsyLA4mzyW3BglCzNLyUD/
sLOrvAjaVTbsGam71u+ac3K5PGqsbC3V2Ta0/bs68njIzcwG7Ey90iB8OdByIH1J7t7u/dIqVMAa
yCEZzuge4mOza08cu6w7B5tXzaawogIs/ET5XO10052RNi2GwDyxJdUzQdWSwvbKdsVCz87Vaszc
AcB8ID8EWQ2QUSpAW2OGdYfGC93c/eIZ9Uy52rF7tZ67UWUU2wzMA5bT9dibyI5mVbS0MZZZvnL1
VMpkm/xep0dlz8IljQU7FdOBxJrQGtRz/kkYZi2PIJTd2KJBaZiZQgxYabXkZpNXOCVRNTaHORZi
zOc3wW++ReGJfAA5yd5qV2tf728NK4Zv1nL4iQ+3kby3MzhIual+YRnOevoloE629a7fS/r16nNP
Q9x0Rv7UxFVymi7o6E2XJ5I4Q98Xr3mfVN1/yqUOS9NcuSX7okHiwTwRJOGXLs6tkNo75In5739y
BLYRs+lb0wRXN+g0OFlHvVH0bR58VRmOX2Fv3o+aUpVwJic5laqeZrLZdgBbAJYQoqoArIk4Owpt
3BjaioKrz80ok0RjY9i0IPufBk52ZrZncKmeMqtGqUlAvUESpftjT4ZNPK5G7f2ovNJWZTkutjHH
FepuVr7zC/vFnBAlzziUlLt+PSAvsVNPwWcDqxsNUd381+HYgNBFsfvheSRgFUM+hQE0UdJtFGbr
9CzEwv3oZrlZCIca7mFX6dQPslp7oZULwjwyuNmgO9p02M2jC2ccKD/kSUG7IxtukUXSc02dbUug
zHrq3zofvw+xLXjRdREfPUssdtAeYKwRpYqDyFwzF+zLR8yS7KOvOAniMPSa4cPMEieTGIz8VJQu
mmhEt6/cXio7sfa2xjoAoLOVDhC6eXcPXezg2tKBhSz/TLX9sltyxJgM2QzcGY1MMel6eHg/HTEr
HKU8fOjcGoWBuw4rKjyW7M15/W720/ib8+3xJnb/iUzrHcgN8a9XCqKAWBa3gnPtSFFNQvbJ5vJT
p8fGC83n9n+hW2ZvSTVKuD480vWkdq3O0daefgdt8wRRMpoGvwRUm24hbPjCKJKKP/gOY7e+YQJq
oTyg3JZvby51GPzlRYJHlXRKRwcn0X6Ahb5we7ii6/yMMfLoDLxiEGY/ds48LSABIElH6ar9RvqL
9/OI7Z3gw00rdvdWYcAQ0BuMYDAPvvLUidkxPTC/DUR5Ikb1eTd9r5wkLEkOTzG84Tjadft33+pv
SGzIcAHEgg1giVo8qWyIH+uMoDnWo07Xj7j3KpyEZHbLnAr5x4dfvecbB71N62f3AtJoZiPTWYKJ
/CapWsh7n3G34HiTTS5GkI3xt7aVBQQDNX9Rrox5jbbh+0cXpkujxInHa7aJbczpTQ3W2rkYaI8P
qteXm6e6Py6G8t4s5WPwIfafsCSbSEpe50N3T+awSOLVtDqF5okZLQKMaBjarFleKDVOT0c6d26B
C9PbtXtUuOI13isuhosUY1+rRPqt1XcDOVSzPGoPV15dksmf3fV7rKgcTQKhmau/hlufVONqvkby
1yB9z+vfjkIplNzBf3uVZNUihw29PYrbOH7XqyzHHX5AHl9W4eeiP5Rnd8XxKhavgF2f8EPFMvBF
oZ6Zv9ijx3IuuyU3SXaR7wzKPaDbGgs4EyJk2xgLdCdjjwsgZrgTRCLiGC+VknsiSA+ipFUmky8I
O95Qt/KXQCyY4EVfVGkaKaneOyV/fxsKcL8Qs3Hhm8pP+Eve3ePXVHGmPiAITsYrO5r4uVjC9kjF
QtzzUwCxu5oPvS50ZyGvRN3sbkn1M92lGCyo0Ui2ecdsnAk0qG+iX/Kw1zs3g95WKB3mX3dYxESY
ky+1G+fGtIfcFi1llYKe8LDR8BQji2vY1utxDeDRBdI694VLt/xeZUse4HSr9hzRA+8PsJHvwYnS
uWqzACU5yVJoQvaSRlqNISk4SckG3f8PDTiL5gErLwFekI7UMg/9vVw6b/WHh3mEtdxVvK3NlD3L
1de26PqqvkLjs+gfIZ3Bs5t2TAyw8iQl3T/6Mo+IQ5fLuCrStiC85mlNkQFYgq9WSmm74XFEEenF
gmCfiH0zAcRM4Jk2pSELEcyurBaH9s306jMgbkxkumu/pymGi5Uuix0HNwjfcm6RcAtD5ZQd8RPR
FVAhcbjZyYJTOoLh7/VkHankXo+xt0Tpss+1twJtbCSe/sK277D2mqFc+je8aNgVh8xNBYuTPkoU
lfBnzjHkB4049xp9/nNHz8+i4Rqnu1By032GDVfJZh/l0Jh1BJFS945iWA8kWhyoK2ZjG/dMRz86
cLIv4U9RG8fXw4+YwS/nzTfPgLgXEPizzL5+JBLPsk7VeYFkEGNSIZuAkpsdqndVzZQeJQOUOG7X
tmxjumN7sKfvClee2rppInuZcAMQ4NDMFDNKsnIG3yppjQBSrJmR2ufvcvIbcQKl/M0cF0RL9e4B
/YLFJ7/8fXbGlqi15/2e9kOFHHZXbUMmZX8VFqh3Summ0zRwl6gdBqSh4Dcqi4sRQYPQNVvDjPQA
rTWITj2pzon3jXj93hFdLWYKI4do18VFG6ElkPFQ774yUql7TDcd5Mc1L2KI6fXT23FrkBXZ1yf6
32hsqilTwbQoLhw3c34jJzAMRhwce+65mu9vYbBXcGkU2ZAb96qxg7f6JDvx+SI6pkVvC4yQr8Ta
CqT+XmhkAs9KYYfnS/W5PolQajO2kLfj8ODmtSGWXrNAZJ1pVtrLBILV4lGRrhuwMuRpgYSkg9BI
dYrOwKc1LY6hW3ZZTRbMNGT9UP6EFJK4rlpvqWvrM/ID5uGiK4UEyeVixVZ3DXPDLseHFJsG840J
LHiOVmvVX0BcRnRTGi4zYB1bUPLyBYxEoQJ2C7yvT+MqQcLIXTmIPy+NlE1DoP7+p/RRuHe0TQO9
Cuo52wdAK/TjWwVBt6iEx3m8mBOYYaeXQ4C5rzbLqQNDXLS5KerQ25E+kwfbSa0aWXGvnNMtOleA
OHXWFWWofXGlC6X07Gjj0IfFwawj5FtTNFNftamedwTNqqMvXdJn3tHyHVpPpa9Z0XW4FVw7STw8
UUNP9zMNQaBE0335ATS0tJkDSGHB/NWDD4N2oxHIPEd1nycaxtQX76e7fm2HoL/JkedOeqnROe5n
GzrCaMBOrOWZ/OTl4gdJB5dTTcSRP8tds0JoqTUh0nKwTnsO8g3G8JOBPsaNkpS66eHpT3Pbv61K
HBtoobKdG2Msi+uz02bQoTX1UZbEK/C+UNbk1EiRl4JC+6ZyqP2x2BAVJxV+xkGkBjqsO1sSK6ND
RM7m6d6ODTf5F57jD2iH/uuDnaj6PWauNzCWSTFPe2hH9Ij3JcrFx6baGDtrOQdd/0qSRWfLFsNq
4qmF+y+wqECNCr66X+IGCf5ux0BMTI4mXpJPb4f6A+PVm0oV3JM1APr6bNVdTCSam7LbXfKghgxU
wDKvPCPtPHN/m5pz5upzFzRQ1Rmfj25QwfVqUQqsxkMW+6VouAOeZ/RX7/bFyvv4g0i93tEVJC7t
divaamru/glgwJrF79vvYGhyTazhxD+ttbf5t8YT4QA7vYi8Mq2H+YTWtfJfj8hZ3idYpLM3W0la
Nm7bQS6ZKLyo+sLHjavMRwc/nKzH6JHizfffrQrDKnnxLjHl3no+NXkHaoK/wpgfUQFcOl0NgOka
pA9EY9r4CWXryw0MRazW8Kmi/+LgJWbaChTjcx5qnykJYnlFEQJkP3dQljw/DxhId8t7Oxa2RMUF
jnVwyW+4RXoIg1Cqdf+Xhx8azX1ziOPUCKhT/skDy9PJO4tEZYs2u2TqAiyYRojYSTcGOmP0Mj0p
YKd8tabpQOwhLw5CCOqIEB2jYZ/ej9bUkGdcsT4916ivuN4TVrtmbyoYc+stiH+IS+aij+O363wN
5avSPVPTTjD/+4WrWaYSLnrZi8WCpNpwFcW8GJnLKMvAkCXRg2OosvSIOfXl9LZoZTLHzznfZiQk
G/NqjWIMjFHCBmf/68uHNuZNGjhLhpIxuU3NMHQYpovM4GBHbaXO4VhKt6vkMuQ+syfsAFQwWPUp
iNW7Lb5LpBr32cVOLkBoukuca3Kr3zIeu6Z0lG0gcO33wYGF8x6CtSaLnhnl0bQbZUVLtDo9VoW8
paxTMcz9wx1/3qCWIMD5dJucbtCcGhh3nw+YdCTibZSnXEWI6AF8kh4ws/sunGCdY1YabmJJK6z4
3KQGx6ntRTNUIBYkDGLXAFwg+ZUUc8S9N37HHcipql1qnRphl8Y2cc8LWkWnPuaFMFRBcAU0oJCn
smpmMuByO5nTLccylaaTVZ575RU2whTWJFhsV3ctx7JaCiQMx0+g9RdDbJvjVao77HzSWJNtr8Er
q+BIhxCMcwnmtBkj7wv4FFZisckCCXD3lVSuPF++8s5n8WTHQI0B0GoDoO4SrY7EFOooY9e2n55O
/JaLvGyYdLVHAa74S3VBUVCk4aghp4QvPCEJ9isAoDuEPkMMvA5FHcSmJ2EXSEz/U/cMpF2w9w/y
mFGaeCq4QnI0sSpMU5fcJjgZUVojgF6Fewb1QHSxtdsc5zNx+bF3UYSYqO6KTFFmUshZwMeTYgU6
LFNc3ajN5+WQVMgFl9nOnOmZ3rirT631amb0JdLFEznye6+qcokKKfseksLoj9EZS04iLSrUmTD4
dWaaOFB4xWK4hDkVz97pdQfoatIAGn3Np7QDIE8nzOzErzRNG9OoO3/SCRWpv9+mtIprPb/CtJNf
gi8v/nNkpO1DdG9QIWUd7zhmhJD/yQrfzSEIFT8UvuRxUfd7O6/+7U0sKrVHLt6w1+RVEG9nAGFR
IDmlAdMHLiaiLDonPlZ8Az2PZBEDQIZSkPUWl8y747drBuigMnPDOMqt+fzVy6BEQL8eQPzwDxCO
6Nr8N9LmgWuoVff1y1EMJvk0C3AiBjRZCTKFN3UqsXdt/PLlRG5pltUN65+KpGPsu8m2AQQWu5Tu
BWoOotn3uPqkLD0P4qa5THqhCAMnT0/xtiWVsq2EaV/yPhQsAtw27VvtRk2ZmC3lAFC/Q5eNkVIG
w3sqzaxu83KtE40/T87mvaib8UjTrD1a28HsBzh2uJuwPcZ6QG1Zgn6BH6A3kOxhmiN6SWRjZaNp
1Wrg3NzPTDEmzMQokjEH1SonOkC3QYVhCWWpNUuDbY9jWSVCrO4uAbbKIJHlKYseN9FSjf9e8m1a
jF/wx+7G/CBvhQoTT/M9zmNI8JBYtarHOVGKOnIsSqx8F1PHM157QBmREDz3SejzQIhyQ7JI/uA+
R7CMqNu5ExxF3JYfq9cpg/XOZosokGP3mpwd6Jec5wAz5hQqNeJTFj7eIsNXUlYrFu5lk8poRLOy
Rg1XKcT1kX9eHN7JLZ6gZGhX2faZ7cHuqi9SJy/dkFyl8aOcQaPpCBCprgoip+nFx2LWEP87KqEW
ZMeUgVzNR9BeWcno4SfwAr6V/NJ4Te+0uICFlvHqCpvKK3AE4BAr8uBk90n617GZ2Cazo3HDdMnL
U4YBAFvfFKd4Cfxzk8aKSgDxD38Ku+OS+LqY630oFDN/QvTcdEZhmNphAyugBN5NCNIf19nXqfNc
W4M/INA1dEMzi8niyshrFhtXTeK2XKMPGfbQpbEkbwsEIoH9ciI+MTByfXzI3u7RqGKlcrXopHUE
fUqwFRFGNW9rNY254YncXRSHi+XedtwVHQnZpn63gmj9iWvABmg44V44nVgWV2+Vab29SSLMKkr2
gJsmN2E6rCtUopS1b9BT4qIAODbdWwQhTPRbt6EgJnkKMCCP5XuA889l3XsNSEcxpRE6GqZo9g+W
GQyr+R8DdHunvPQZeOV5SKX2+OUdMB0te7HMN1g6adYgxODlqCA3Um2hH7AhK0sLu0gTq0MKVEos
Y3lUVEysWWEhHIBAPWi7iSgDLdvFIyRC9ahZeM/7n2R6SpvhkCHctlH6FsongcRQbdh5/P/a60tB
t5DL3eRi7IK42NE0EVDtlj5nzLfYNrL/BB+2TzSWY3QOvLSFg9TYo5/vPAHmV9BJZ7gM5+RSq3FH
N6AjAI2q92+wUyaz4VbMDDLHyyzK5T1QYmOzEln39zR2ZsFCybduX2MjtPshYNR1FYIWBjSSWuYP
kKXKrydB/qsdZe2FjAaF/ygx78h+C9gPGXlsIp6CxsXp1pWNYLNswBb4wRCnUI0LAHgg7uu9SRVK
2dtul4ImXkW6z4Ud2Ur4ODTpRnxihxiB64+dDToGudNfQ+rHpQsYPAtHYamVJTEl5g5XBVnRdDLc
Wwb02fGB6OyXxZyrdlsk0tTWPGyX7ZNcN6RVzdkKdO3a15mbR8FYM420VhFPGpWwloDj3C2pX40i
kAvhI1OzF8snd7nkuihTp9eK/PGTj7J4gIsc5v3LSaKMx/qdd8XoSJtwPmh3gM0KJ49nO9sdQSHc
+ESWYZWYMleDpxzUL3uu8m55u4hG0gBgH5lpTuJY+7SOq+GEL0iPB2xK2krEOxTJUan4NAEars1T
miDeBGZcV20SQS20QyisGBg/KZLP7SorjjwZQdQ1xjTHRa+JW7CzSnSYyI+6YuoRwjNvwz0UXRSR
kQX6vy8dJCf+PFf5jfV39UVM85g80p8GN+5u/q4XYrwCm74sESnwEuKQMFFDOkkq+9Ff1CwTdPO2
ZcGXTWCpfBuKkjzTsexl/ig3n88LoJg+tYKuEKyZINdBOzzUhKR8V3/n3SEddspzbtohd8JNK8Lj
5nmLteigsM5W2MkH9Ww5yLc398vxdheMQqJhOJ++8WaPgv0yAwEY6lSj+1S93KPILKuLLE6j48FG
uDd79st+MxJ8SKPydwYm85R47Or+tNpnUdIxxOv2JMLCiNfOuIWHgw0bzR8sB/6Cdc7qF7hm0SL1
9OGL83f9J25ZV0i9Fmaq4cJ8hTorGRTuRD7fpo40ZukosI858sDEuVn4TEOyg2olxjTKp6pV2za4
MN0/uQIQwVBWF1IRsSwokEyN6Qfq+FirC+4Fl8Kjfkm2O5Y82wIahcgImrAppaiz4RTuKS8IcQNe
qaxdbrDAqL428VGrBNchwjU/eC1IBesLHH9gQIvsigepecqePppJLSQPZEKVIvLStb2hM29qaf8F
u4qDttylqoqW96pm5+QrnCO1hOqCwZ71iOTeRoZ9u0b5xVt/1rXASfPxE7sPMI9ScnwE4kFLRi7w
bR5DkwNZBCoFBR6CHp2jJTsk3iq5GSdpkx3e/3pfbT9vDnkpzhRRQMkUpfJNLC2hYJNm+QumFQjF
F1zKm01vC2RdO9wfTeO2PBue6t04pgmDmskG1XFFz81AXivkG/iQ2ThsCFvU3COtNf3JbAz1QqKc
nd34iEwmYBV+ntEi+57Z2vQH5W3HfeSyM96LytWtrdHWhIgZRdSQJuOuplne4sEyCc/FVBkKmFKZ
sWsdJEvvmzkxCMgGPpd7Cgi/Cqj+mY8IEjDA8y9+4Lb9xGxY+Aj45LaDNSKBYuAOzzodO/bMJuQL
CZ+U3Tgp4eptUTX9Z4wwv08NuO9ACl2otLW6s+Jx9VbCjgsBFMZA7F3FRrrF45KKOyx7n54fE6zT
faAezPfSg7IEJXtT4SW12QU2uSbfUPKydlflri5UYodvO6rnipSz/zEFqgbdbz5QM/DhggmbuHPf
HCDAcMwzI9R3c8zVHybccISyTDrrVeqlDZ8LfWYeonNh5LuezR/HBlaxEBI/4g1Qc4DcpU8P5at6
dHdNpQGuBH4OJC2KLE1WXEs/2SqcvPIRXY25lK53Fch5Li8aAoJHNXM9ODbKCTFa/ci7I/YysUna
7gpGiYI0dqzAwBUD2Gy386j+aeJWbJv50rEHYU5i7PzUsIRIu6KKou/qs898OS33F4Jau0DHw+Bu
fTek5VMIYVNpNZ5XiJsGJb2xSd4k1xDVSk0Sh+q1T0X3reYt9Q/VQhXeLFfvljBbMociTHZKDDXP
T1LyHEXLyVByAFaJrxdPU94CRHrxn38EMFbjYFJ1YST32wznwHF2vj35UNEfRuRhIDnl2Gqe4QHF
2qoLiWOk8CrIPtDxN7Dnd6hcTZW4z4EMlRX2CHGFPEQ7ZkiLw+CUwSwDUF/r6dhBeGVSfniZMwzw
PsSrqdf9FgPpr/wu8ODO6cAkbJeLMhsFlMh25UWY9ETawkwH1FuF1PqSUT7TyGaOT7q7nV0cMD+q
UjlUqxpkxKtiNWIRopBebIyGmpzsBPZJ/xBdFqyWXpRYkuBDrpFXJrXmzZqvjxFSr+q9QWshOis4
OIA3R5fKt6eZqVsA2mH+prWls/cvpugi1c64hoegorF8R92ug3MEq7FFtkIAWTz/+PPm4eoIqiCF
X0OFNNyd0uY4XmhMPDtWl4M/hC5iFHgGWgbGPom3W3FTkspPzLKWpdgPDKxELCWzZb4EB/Md2Xdu
axrYjMyehh1kjFIIWVt+SIfD33Vra69HGqvzGSYu4/ZCz9gPXAoyUJPtCziBJLGt23/G1rUmTIVi
SDEYrhHaFOWklXaMErrYt8RX+JagPtl37lL9gJ9airFLUOguwdnipt3Bn7cUfOyaCVqmUj/c5Jwh
1wsu0IFiVE9LvQO68u8FCOg/CMoUNBDOFR6dpWLxud7VxvOVOoZczrGTZLySJ4r1fAxhnvSiw+Zj
vBmRj3nY/T2qAmt/OBEU0umNyNeOWBs2koKidI/rrLw7gdLLkQAwcX05LAhZBSX19qsjBN/O1q72
6csoYd51xzcmIBnGT1nTVubjb4WZZgd7k2p82Wg7f9Us/gvv/XYcPjG7kuawndEXydp9WP110OYG
n+13u/xyugk3fOPoUzdUNOihZ77Z4tF3fwLxsGoSz2IXeqokeYHFAmlTNemu+Qnj7UlPLCBXXdox
qG+4zu+GWYgQqKSYPbfzMg2ItGNQXdpUMc+/I1W26pBuNexmoFyK+eY0t/HytZwzzYGftbzt1UCM
mi+IbuM8am2b1M8YueJ0L9F4Y0EP7NFFnLB+Dhi/d3ALPIEeqjcJZdmrJjwGXVSE0ONKFq7D/t4J
+pWKtVUSH4azsFvq11rAVFlD/Pg4L5qG9l7owXeQSEqL8i87hVBCK6SgvSAsU1HJQD08B1aYVsUl
/9NO+Chq6H/ZP2MnHFuudVLQOtlRXs037t4wAinKo5DDTH00Wy+chAdFWOfrHbaFrWLG7nJDqIPU
CYw7ZqUtQoHl/+9R0MlXC+iWEosD7kIZnWNxQMwHksyL53htPaol7JCVIIR5y+2fV/0i4mqY+Naj
zX4DSXa9cOKm7GFABh0m+8NBJxUokgZ/FeL8wcDCPsBkoL+LJyE8wqXzPCm5JJrPySzV2ax5b42w
HuKn+9QA/yO/Azf/GoYTR0zSXtzzahBPkHsYJKXiPqioek1pHOSqJqqJaF8a/ZqILVnSVbw6FrH6
bAId+35dAb/04OlBLzEp9KhEhXAYomozNfvouEgReIH3AlmkgiNU4XNBZohdu4rskCNyJegyyI4K
djV6ozGcgiFlsP3QCAd5wtBUzu8zu1DuYewIYYq5OPFdDcNcOJRjiEeyVyShvu6JtTSq8S4Y7uvW
q1KlxnQts9VknI49k/6KV4oMOS70tpAQ67KR2qXEmtArBIEuUxG2a5wXSK6cf+thLA4xJCDK0kGM
nywSlunVVTAUblG8yaCeTqGD70+R+Gtv2nqeiPCmw8BBRDSwrBzOIqBn/uCHw4Ra++2sYpa2OZvO
Q2B0ggAHml73Pkr4M0paMBnpL+05qhYPE6Iu19QvNLskqEuBrZH/61AtRiQbIsq81p0X6E6PUCp/
oiihXJNNHPH7/APYKYIBK7L7oQj9jMlWOy+d9PZlODL9Qy3LgoRCwi1aq8vVSrjUTPy0MAfo+NGm
bDyl9W2QzJoFPwtLABerFsjz2c2JXf0CWjqbqmcpsLfthEwqJicsmwnIwvyqrbH628paGIXd8V58
EOZZeuoNpm7fRM2W9fUe3EX6Zvi0dJXlZH+bhYwpi5ofm1k+h8BUGkMl6fbt7ssCa/0Z7JkAVeay
j6KwhoYDRFoBfuewPOE7s3Z9KU521OukvDW1FqcD8rHWCv9Cu6KDlL/81K23GCe6ONI35g3LvOTp
NKGjV+s/igi5v8kagPVMtVv9u7sw5cszV8xgeKFRFxWChKGINp0amu6BPvdu1fERZo6lVldPZVRM
pFCdgWMb3jlVXOwQUz0KPKOmbDtTkDyy5UCwpI+6gSaVRT0M1fMoVPEYLq/mafAAa8nKCc+vc9zT
oJDZeYAdQtSKvWW0DSvWnn0Qri/zYfqhvS0MQkgatTexNohIyQ+zz7FXwbNvc/kvDc9GONfb7Dky
+f0Q09bI7L73eFUWwqdH7wi2ua2dSrDV7k72si/ekh+SlxjTXVzM2zPuKAlWDYzD9qceD1935HEy
6hnT3bFQlKuJyHqOaH+AAU6L8v6unWSB7NQk4WQ4f5hwg0LwGcJGLm/LLi5V+a/e3Pw8cQD4J+Lw
4fbPk980CRZQOvVGx5nnPs7kYX8UJGSg24uFLzZwnX74//5EQfYUzZFWNnGTSrMA681Z/WRi1uBl
KJhZZGq0RXAE8YJJCVpnTc/uueFeDqV2lQDIILq83UYgCV087l8Py+lD8byPmizNM4imo2/+nPKx
ekYkM0DDYgPNWzCrbwj/ZqPcU422Eqsoj+S5r5UlivEE8sqVFeVrbALnuT2i/5xnAbMQlvXwaXja
iT3UihybkuX8E5ahcIFMrI10d/oleymAqHZB1T4fo2R19pC7tDCIX47/XMQYbmX90For4wjhv2Li
fn/b8rdY6J/AZHl83rZ1/cK/Tuu/7ZY0aELKtKjLcxihULPInHjm0gx/TYGanPpYZEhxKbR30gup
JWS6sqWbeXRY5/B9FBjvy7EVCTJxBS1teq1j1UQ6k6cIibmPrFOEvY/gFKTK5RJBaQHKE1BvvOKS
ibFdfPM1UfFGYy23QgsDr2whpiUyl/uf+/Yb6rL1LVDqxgUJ919FFQr0AarNcRM1I6kna3N2ifMm
mqoecR7JqrR2Pid/eZrIwdLQPwwCtCVFZRByheP0fQu8ci+b/ug7nviNTWtCN71iTO1PDFpdtuOD
z4peNu+VyWi+ohIiVhAuQdPuQYsdZvBb6uVtFxM5pXCg+sUyM4yPKyKIKD0Drk1kaHD+ggtaxbv6
U068rXdMDUDW1PzyIPQU9ZtEWMGLq+VhVGVUq/OFFMxwPb6Wf7UQ6NXAYmln95LluDR86S9fFuEF
HB3bXO4jIQGTmCadx37mFG8eZOZGFGbOWSvQl7ahsdNoRq1YwWAUE09DG+cnK4CFOJ7ugwxJ152h
pFQf3tVSisGlwZQOhNVOXdQefaR5v/qcVJ6mUZJrcLJB6kQ5KqQ3Oof7Z83hz3qaMTYgduG9DO6B
etDKhcIjL7TubFBRt0JETchJwDD6GDmlw/IiVIbxa2wALrcM/S+DUThQWqedGoTwMFnkeKVTji/j
LLwh6++fJIhsGnyDJ4k39h0vRth5NboXBD7qIXxEITmCBe/tuRSW7swmVyW9wYfme+tfTYQXhNIZ
JZ5p8YJ6fU1Zxa1Xd5mX5wk/nRfwhvepVDLTbSRXAqMCrFOC4KiXIiJrQjr4gt5FUhVmlg1Ya1LR
i08WP+Cp6P8Placgp/wy7/hvPzSXzdmbVD8d8S7Yvzem+jcTeGUnRnxrEz5c9F9BXOKltTjysM8P
G9nTsL9UKfBZX+n8rOEeIsLPAUet3klt4onUwvK8aSlaoA8wC2S2pgeFp4uAxcK8HXPQMjTOZuxK
Hxq5yC8f14dEYMrLMj2TrJ30Jj/FaE+5R9Fx3Cd94q3qdgrkQyW8p3ABS4jghKCFW2FUxvl6t2+h
MCkDludLHbmoQwAc8OjE7oq4PNXGxk5Pmvo/V1BZp0vX3AgU8j36X4I5MptDaWLKXMlGYwtnXvz7
2YWRsRQG2z0Bk5TSBnHnYtZdpGSb9na1sWD4oWfl8OAiTJNlD6sa+zaPnj+jkZQfEPvVhB674V4M
av/uPeNn+owgtj1gpHZXX3j0wuY3/3Vv7iUJP6QASpWYZif4ooeiKjCl/4T7e6hE1M1fSNuPAHax
KCNGiJoGfk4snaxRsaQ6Qu+Un1r/iHvQ+8CmRCK9cj+LdLBgm19MrVjyy0NuWvcKVs2fTYKTP9UO
NU9ZRAjJ+0WKJwjjql3R4BramP6DnTBQOnKZjDK3SHkyO/+b+h0SIrtVsVG51WdBCQ2v/vBnkk4B
BENDBTNP7I7RyD7LabJEI15xLDUWN9z7GlzQP+01fParOaXWONSkQjj3NrAwTBMzfKMdSjpcvkEu
XYvr+n7T9+SOVtM3NdnhZW7+yMhGvB2Ld5eABSG1mkw8+10DAyHkgPnDbJjrq9ST/cc47BYFN3s/
ZO4Gg/EViSSjwR9TATUhTY5ysuTeYSiSwSZVXKI4AV7f2SrgfDt6RMsgg+OEeV5Yar7dhizJOJ7M
rxMAUsinyxf+Za3Fm/GD6ZXFOm5lUIUGt5zNy1rJFqx2f+GUau16ID2eJ5FHMWWofSzUVIhah6Ik
sKNyBb2S7WkLtVPbeOjNRSEd8w/Y8zkyyl6UV0/E3LgRy6wAJGTtIPg9nTLH/9MtwHt/wqNffTsO
ENxtZwlrmFeguvApy6D7Ye5nJmQFYNti92cSWDc3/2+kMZ6c9EGxqazaB7wkm/qmhg8Dr8Ap2Z6C
2e2pK+rLME812yCcWnv4gzqgY5YdPEOtkebIBTK7gB4phNi2qNHwO2K5AeWNZ2NNH5INmb75ef2v
xVxIiRhIqW0b2hgYFzqX6W07La2sWr2Gish4PHaeYMsVPzhsSIhRn66pUREOVAXPVrejhvbjwQi3
GNXbPHds63Vrwf70pI+JXHHoQ11z3qA054UX9k/SzUXTT1EQabb6JlXQI8sxLvVzlVLUB0Fo2SSk
qSHXlOh1nJUIJIyVE/I5l1O/dzC4frML4sBKMPZPhjEGxe6/YJRsEj9/w0LXEfyp76TRQ7k70XKf
GYdfOXJtbnaBJyMU9dzsqaeN2Q3/6FtOgKtLeggOXJYVdMTUbbqCUplU1gIBuwWEAaMXG5cEKzFd
ivNGQX7yK4fDb5gclIDHfrOHszjcPmywhsPFksbGkVKwmIIN6B0qpOG3rzYNyMH0kflwM7rO06vp
m9of0QGgy8FphmTO/8vPJTCNJ3N/jxr1dpRdgkh0z752/vx4VoVnn6FwUmV2j5L0XPNW0K3L1cy8
0XeF+3D1iZ5pMfotPJEZaFirGOGIfmV3WpBVC2me3zgMMMjbweR3/sEgvjSyiwe2kaAPjNtXoa7b
sWlqrGO2lNAOIq55N9YzJsm4iQioYJWjuQwVdvHS7SQkGyKL4B5552rjkPZ4tDfTkrMHhrl1CCfg
uln22ajCalupWU2Q5qqlMhOjnb89RQlibb1oHc0E4K8F3nn3lKo6a76t9zSv474NnLEFw0nOOCAe
EmYgmifZpf4l+B93kRtv3k4iAuXhjIt/NHsY3KoU4DBezeV4f2goE+lpTv494bmIHfYhGrSmy0KB
/ANftsKO41NPqrJsMkBETVg3BdXWuK/kG3bP08yrhGi1dmNsqKKw9AbuaYHTYqmzfDs3hIkcMuAO
RtoYvG12JEv542L0ljO6fMDzVWMAJIJ5z+bs0aPVQr8pJyVfNvAESLLZtawt1DhLFXNBxnb99eLt
oPaiFMOkUL27z/DOMa5HupW1n2moCRWcL8mOq6EdFfNftOdFyup6NMKSG+gxe9xUVoGp8/axrwXe
47jINVDubDmSqbYN9UPPwwQAM7jsDRrVERqmLsMmoRMkqt32UejixC+y8+z3xJCjIkb0wJr1CGLS
cb6gFnGPvtK+XMe25vhT4yCwM+WpZGuckK7L/dweuAdiNUkljFsC98amfZ+g/0OYnKO9Y0MZwPgn
6anyEM2jKHEKKvkBVnkQAMKtUKHsK9L+AlXXwF0ogdbRQPfVWRrV/I3PSSykzpSsR5P+2k0Q9Iq5
XAg8yShxpD5kCNhmfVQRGV8KIV/VEndq9xMDnB6LqPtF+EwL5XsfZRyubHh5a2vaXyGDP8ORSMTr
i6cjky/2NgGlV9cB5N7wjHMNVngejmPouKhSAyyLL2n5nKjZhSUs194CuWdPobEpcZFuXUZpYTRV
1eCkwXnhNZEw+ClK0Zd+kkLmy7n97BT+gt3Y3E3g62np62f05tPbTMVT0wrsaQtvdRQeqaQf5I9u
qgCCkhUeJXKw+5Xeqj6puRUlIhQFszY/7KqAHFhGwrCg5jaakHyMavUqM/LTKbmR1Hw95LWpK5XK
QgLBk2FEBLpfr7TKegcvj7v1q/r0e0kS5gLu3RyboHNfgEeYFbSjeuDLIWUxiXf1X2XDWzX1sqEM
fRepIlFQgmIGot9PcJrs+x62G2maZ6ME5QAoQ/ANp/+8N4id60qvQYzPFB9CB4ucgTrSyK4/ef+E
DYzNZ7KTBlGtRGJYLSPx/G6ySOs920u5iMvh8Wk9Gz6vlpXmSXMKL+EdT4fdeUJ4TZ77E5aV/J2N
HmgLU2irjKrgpXyYSB3JrM+GVeviRvYPKAhOEAUrKo7Ypt4irbZHT/8dT7qUm11iclfy9QCWWMUB
t5aEludMcQLsoTrTE3hWNl/2p0LIXtVwvtmUhoBO/PI9syeVfiYiIisauPtt+fUr00Ly7LijWkKJ
2EK7JJTJL+E7MJJakOOqlCVsxXFjLfNz6Kc/xvd9DafRcruHRG5P50115eN6E1n0Pb4BXQzKPsXr
qTl+Dac+tVN0nxwYiItIQflzsy6mdh6pd+nUDjR4dQSuL4DDLVbRKExMrzQwRPb+ebZCPw18e3T9
6S5sjvQMwVcmGh8FPgKjjJAktAIoMpXRTlwieJ9Ewtnk5mQtfK9bbKc27os2uUGQ0ebc+i2N3+kc
/452V6qAfV8NbYLxxPmgSiI4KUHoBhLoyDGkIOCD3dIg8DgBLj0e9E8bwlX0AsTKpS2x269EFy+9
MlnfYQH4wnneuMGbLLHuG5yZXfMwshDIV8B+GXM++Auosds83+SOlR8mlmQQ1PP22dlFzHlP0xqf
vqi8PDDNl1nSNaAMkwGc25xOjg8QCiBwiUdaphRXgEUmS7lvavNqdezEY8qqxUoAuPr5R45xHbF1
A98OGK/03Sf1MaZh8ga/HQXvjlZeh9upHJttaoamRL52hzXnLNUj5ptgh3yuUYhUNCrvtgcYtdC2
kjdkwNgTQvWmyDyjofZRIubHXiZeETKJNuYZq0Zct+x2P37Ue9r+/aCgOT3uhSFbyQAsT1XXXYhD
XRrhIyyrPxJh1TDt4O7v8HsFXNuF/bZDGxml+vn7Yb7msaRXMDgKpUONTKbMNNjCTB9OI9kBDYYq
tUoiREZBxz5bGkT28/44WlUot4Z1f7mg5fcpSlG/BCLC4Yr8pQKqSUtFPcSSco0agcnyuXOm4WKP
445bhBSTUzy2NR67siyyd5YVa/fF7X/cjAUsyNg7844cIsk7Hcs/12epPeHmatQc74f2rkDZ9JrF
QGc5LTU/E5nYoolkogjOT+NH1WHKR7PDaM6H3QYA3RzLq9/HDv3MJXosck86e9X7sdkU6D4G03EL
Zo5232Zhijgtb8AyR/pgtkBZpzcBL/xwU45JMllKgoUgJeVaa8Cs/nEVMR27tNyK50rrwKz4ulqV
Od0zHD4AVSTp7xtS2hkGU0qyjT6QMIRc8ebpnd22bMFVTcP7GiIhVicwMf+4xGG9AVWhESoaCGJf
4tImXrsTgAx0ECWDJGW9Y74VhjWNJhQlCWhmiDljErIFd31Ugd18ZIAKSZ2b95av6Lh78jr3y83y
mXQq0K0MB+ddeeOWzuX5gbEKV94WfOXVfwVSCC4QYoB63jQeOssA5z6qf2KXb7jgOk+AUn+XWzWI
7jfJdEIiEi3MADB0ce4Wbrtae4/TwxtBLqjKPKSassh1qRZ/Assa30AgaAy1eJvGP+1tQw5y14TG
/YMtFobyGxxIjbowwmSqdN7zzhav9+aNDSw41IGXhpO+Ck2EO3Iq3R7EHobfNkSLrgHPP1gC5zXE
tGrrbdKZhtuEfrswyyPP2q045u8RTk4agUSt07wnDN9jbeTzdd8lCvQ/WgeUDdFBAuaIAbpqMjgN
/5usW6YiTDQ7ZH4bKyIlg54ING6mVid7unVGrvXMw4UZh40oBi4830A2e5RfcH4GXjJrOOgH8ssl
eXKQVYBjsrsKzLZ5Y9jGvniIOXWOj8dcfErWNslPInho9DfXSp57sYHqtKPpwyngfK5nkO8M1JYC
+qo7bugy1ulcY8qJ88FyDXmJSE9ua0WtWWEp/EWcVKJhKRfwfSV1tFb5PSV/0oOS9U+t59KnA8HJ
4NzztG9wZXNC3dwmhMjH6lC8DEvDXoPFOPoZB0MIyD7r2+WD2xxBPaq1dNS3VAcpOLVsGgo8He9i
2ApWBK4d6YVQI4M8UDEJzXt4yYxyeKRJJl9ZSDPqvPIwVm+ovuOIT9a4jN450mTSInxkpIATWnPX
7QnGXadjcoCwAaNPCtIg873HXGwWsUNwJSBWfHSRqoPcH168Sg71TmBBDGDAVn/9/7lWnADUI2vl
Q+oBw9jPwHOtD/CwsNvuZ21l5kSOSDQYtis4zcUH5AZaFNDWlu8KBQzKGrNzHMyuGJmD+ftNj6pK
StVzCoPX9d8zHlyjROGBIeEwO8/WUfJB732DjcKYHzpa+swVtqcIwAvg81wFEkPfK2Sw+MSdVOz/
HVhrfWM4z4D5og0PrHuWIZYvnUzgjA/0dC/ap8G8UuR6x8xS7F48+Fi89N0OIgO4Sp9EI3QlKOmw
nseIulmaghzcbJMwCmR81OvABs3ADUsJqRme8ctHYeYd1Ezs+eJg4jMCnVOpEyH/YVQ4bNiMjznz
embtVtwWZn00H9JvQw+M+qsYnbp8Yv3cItBbs2ko/fdakkJd/Kn+9Yd8CAN23CY0mN6+2DkWsX18
mA61DJfkpLuN+4av6zcHvTmkkC9NYzWfApo8+JXO9pfUMwxjJQa00mlEfQfReL36zhuPySXtHgfy
/LFxahOWQh3C8x/h6P/4EmOiFH2XlCAWGnU0hAEhBo1aG8TmKS752rERinj0+tSRiJEwkH51/Ebi
z8amUHmuEEKfcbYCM2K2C/MMSqBSp2N//xSCu9OVGQAh7VIIEXEHQ/WQjk66a/i/P4wu52j8VTlb
vEz+9oU6DB3c3y87KeKyD+Rwfwr2xa35ZEJzO2fjNBvBaIXAMGNdHWPMAP19CV3bOaE663Z/6Y93
ih45edvBxXZsVHayGjeITnSvTzJRs8UTuT2AYjUhfBhBtFTNP/mVFgjvBUH+TkIQsofNf8JLZEsa
OmTFUf0L3DHp7lA093YNBBDfdnvUrgm330Pm9kXF8/rBKtcZ1QNtFIYebMoI33hA1lHc1xm3G1y/
ggrLkglqJ4qg5lJ8fLlW3vhDulzwQps19XD7nG3YCFcFCTZGWGm2rUCALDZ2aaGSBDXPiRfQSpw+
2INzt7UctopDlaVaVapuJ/8UGYJm0kbn08aVf8jlWGNg0AyJuSK6NxB8xo3GDM+czS/MCS7+Lh/M
Icv4GtpoDR4XoOYwJTdHYq5g0aptqsFVwpc8ixwK4jGkWn9Mdl9zlykmx0J0vRD050cO+2jxqm6Y
lcav+Spr4LcWEnYUAJCHYTfPBvrJ7SKY+cWPuKg0i0DSKeCsu6lbOCOIc2ouLH+s7RaP96edWZW5
oFsE1SYEjDXOwvrQLK+CjZOTFDobw/hnKYR4JnpFwbYgWCNBCt4ymDdFB6QFwULtY4SznDRkXuw5
0DvYpZfSOjzzLpiCRbP/9dgf2+97xPJEi9bdT7ujrVFElw54kzKMVYXCAuivoHjGTMNRqPvQxRVX
JzAXDTV+icPP5dnqzAjV3A3K6DXbMX8mAdwVG9tvMxiemZLfZSmhUHJLmuM8gMEI19lQMrLiuzu1
/71oGIOjtUw7QFLo+CSRcRMuhDtHfFFcVayyk4LdCLn/DFcHBL4++qiKyFrbIbtBnih67pOs2qL8
oqnyrkWMuRce0R6F3hnOOphOIyLHsk/T6kRmIALHZz+4E+Yk5LfAGkFG6SFT+nt6lZBOB0tCxKb1
0R1A29+oJlNZZIHoq9H8f9kgERBUiME2xt1e7sgiTy6pQw+lUhM/nQL/DQDJvtTCsHmK5CODKJEA
Ug1o0OgTrtc34r6sGHbfVSn2aBtoyMhumc854LIMIl4sY6vaMkrkWZnlQu9B66CEBCVpi9FcQfPm
+IZNreWJXWd95e6nGQroP3bUOhULmcOcryliDeJdewgjGjzowcK/rFmFhwMMMFpAtCqPC+QQA2A4
okA2dcjMj8sdm6Vk0pEMV4oM8vrMOrCIl1BornGO5LBMNtRRXqc7+hD8NCUSpPalwQAG8tEQPRUv
72xAQtarxNSlm7h/lawTsLf9fyF+NjPX/Cg+aaW/RPG4/61FFAEx8aYxeJiwPvgF27Q2qh56QyVu
S56+ShJ9v97B2VDz8uoNyqeuyrFrC4c4hVaZqnjpoSansZQtyDrMnctxcR+Ue7rRezoCpwISMpKD
wz3t0ana8fOPtmnh7fOIC21tKoQ6sdlpiJGuPsJmDzDvR9L2tUwIIjNScUEw3zYahYUNWRo/IWmY
RmvG8YHMpT0f2l/YciZOFHX/8Aa7GCMi0yIR4+RzLXjGWEMeCEnG3RfLMN4ZNw0Zicd3qsuUhyGy
Y59XAP7ezYbKCdP6OrqGCae087tyvHRMuipLKCslbFzlXEtRJhJT+q/l9jybdFOuR6ehKfxRZkF+
xnZhK34wq60aZczvpUHk1Vrzto6WVT2Rp50kL1kXQ//Wwv602LajTYwSQdMzRK7ZVrkdbKor33jv
svBSWSVL85aL/znFbPMUMzkS8YJoNVnDKgQOi5J4QnV2hH6qReh83xaAwh87LH4ZS0LsEoWx6+e3
m+PRyrBoBuCnFgUx8gnt3YnCnYwq1Zwq+f8BBKiJm1ofC9Y4Fs7Ou0HvEgY/ia9sY1DLFxjBdYJH
EuinI7cI4lzVsHkDFsGRskdnGsrjnsjF5LIlO7SVu1VVHvpzvzhK8czWu4WpXfFOGPWDI1uJs0UZ
bNZHUe8jFFIzO2tztezx4jDof8YPYfbv/WzQ+NlqZtkoGpoMPN4GLbbHgFH9Y9/t24CdCPrboaBp
11xbCERoE7fRLl045MAR2TeZ241PcRPo6H5nNJQELbx5aXZpnd25ISHWziAp0/uuooytIxKrQLIE
qOQ6qV1T/TVfqdSs97NRUhggx+Aruaraad0gPAvLMutHrx6dOmoB9bHjOW4DSmQqddZ4dFY60k9Z
eMUl68ZrRx2wawZc05d5ZeE0oIeBT9fM0LQcVPQH/w+cWz9LuX+cilxbSNmOpVNYWC2rW9WG+dWy
8tqYVNWvCSFOf9ItXrvEijJLroSIt4lq+e7+AVmTGSAlzS2naf3UDnqll1PqMiIic3wcN9QniNiX
GURJLff5jgKR+DF3DHWzLpeIDW45MqYnvJo3/a6w7TaFn9sOFs2FOsg40G1GB6RKtq9NqZF8E9X9
XTLYuUu7yFRqEyfJ8TzlPCbxs+r0lMx1+5Hq0y1A5Xktq4vfKKG/4h+PLjdcyCPpdvWtWl1tIFJd
R9YHCWCVDAXv+ZHDOcQ9Arm6U4oM+siY3lzy9QmCjmWoclGSTToAsVfQQZr+3Zj6PqtoGaIs6Fpj
KLCEQoRl0/WPJMo4G9UMVq1Yp9hjB6lah6mbacUtLEPkCK4xG8GARqeqcszwUoDlQ+W8QHVH7CML
X47/Auegxh8kuWK6apBnEhFADsDlZE0QNNDqII5lvyofXYFhGNfPn4GU1qrgaicgQebqigzHkCQJ
0gSBbcjhlrasMzbn0hVycCG2UqvI+e2wSey41qAq3MH9gOObBRKT2x/t4uDp8M8koPPuNDbEB5Y8
41pe1rRjiepzLmccyrefgq4iFTpZHiVu3pPOGIGYu9Bvo9JDORysrAicN6IwLZ4dXEOBWxyST4L3
5vU/3WOFPsh7CQVEZLnYdfJP4bKOunxT1nU7o6y+PjtzOaxm2jp3jjSd2u6OycBZA+9NOOglhn0/
9J6/buHAcrpZsGY42toRBIOA4toMI04OONvXo+GcstCCHpPd7LIaM/iHfyidZZssQwgNZFBTQ2BN
z16O9/iAfcIRvAnJhYRQx9mBdX51rAdT9PhIceDpgvU77MPRaUmtxhOzmON7FLdTHfWBJQYkBBG4
w8H/W1eawE/1dSaz+Iokerg4VcIl8SVWQysVfIfYUyVgG7PHvm0wDzL3Bbf0JOh3FU9+u2bGncqs
02EsSDFDOfiIJfHnjMk5rfO8CimZDkwsy5PZ9wWAn5K3dD9dBxoopnZDCZa4KpvKoOQHt4VmtxSZ
3b4OjzugALSI7CQiloqtSJOY/sjMqVQ3twcl5o/LjSWuAGIlS3WTOs1RRpByaJWeq1jetDpUkl1/
g99iiQ5S8Ojs8boLmcgbvuLWOH0w5zqrUw0fuwzCa8NKUacl5qJVNIaOPgtFyYaeabRyDrz+RpQ2
sDLtIpBtXMV98h7FbDnvlkdSiF5tWuswVVEjyXFklLsDjE+ZOmeuCEQQbR7sLGcRq7odG0Ow7n9N
UE2omo/6AnrP/PEJ461WuR0krOHDcBnLIuWIgHM8/OCm8qGLzD+TnktR6i31vMrspIl+pfy1DC5i
1C88h3mF06i7r0+hWbh/br2BPwRaV0enY1rfh3VJfFK9+ftbFy3vPUUX49bOe7SiwMS361YJ/j6R
CvJgfMUT5u9kv1rnDww+OTXwjkdWtsr4qaCFfJqT9N1a3I6Ea2iUMkAjZ5YUgQEHbszA0vaJa8Q1
6QIZDWI9h94WjKqQLRnZIJQp9oELeYY7SgcScASpOVRZOT4mseErrfysLqNOeQfVZhcr+QPq2QPs
3muL8ilsvTnBHJ3BnWWWcKQJOhIdINt1zQS2ZPPHaCVIh6HrY3Ipu9M6JXrG0Yy+Wlzh+Io4n77d
y1WagB7UWsBAV+mp7q4NuYqxH2rD9qS7icI2Hb67TucyEXbXJP4oEGpVmaOv5IaXZ30bgV2ofnKI
206zLnPXVvrErpbpa3DKBh7UKH2Wh6PfdKOGJhKPbGzAzrFBPaQ45kj12XLBt8BhG59+0sd9mEHS
kFNPtUJ+uPGHQLHKUyMNuOoCk0YTWOjIpYyRwpdSxWCk3kdT2URALzsMX9NmQYimpxzaOBlHqBc3
sTulDKWNjbK0BtGrHdSkW7pTwAW0oejprai+6StKE9QOghyZTWlfUWcv4Q5nrzD1qX8fJTjt8gGY
47cVy2/VKkIvD6MUwGC0fUfKDwDysQeS6nlo7wQ2cRPzXKvnRQTZiJ7szkBXvMBls6feethsRMhN
rkBk4KNfU3ZWQtVUSN+BdswpzqmwfFsbu8LEKZe5ecH+qK2ulTxoQFi9D0vOQ42Iz3ecsiXn0MBk
GJxLg0ikCQ62zkoqbcXN17hYNGPV8LIYjFzGI4Sny2iUMd6400u4nA+u/Pqf8J4UYmYgC2ZjiGrG
kr1r0kQFpmioCXTNFmrpvLDMpt20Bfz7yCnFqJ6GE9tDJ1h/aQ6khGNEQopLkLGNpMPzLoq3De/i
3AiQGLkzkeQgKdrhQcu79YWQaE61U9qEWG21EsW/Lba4mah2aWQ3RlcnRJkM6A95CtEZ1OcErz4u
Fw2TLxHxR5yQyG8j7N+1VTPcNuV8egMuv4JLZ72RL5anZwTsJXclaYUOTM1z6Vd2hEED2SH4Fjjk
JsntFbnAIjrU3gz7Y6subYGfGoQsVtYwUaZ92fJsU+pZzSD4vclPOgIBseoiIva00uQzWG38fEwb
BtxV4t+FQ/dbYPJJK+ZqmkCjPFts+GJvpb6kuzEi9gB1CUQemR2jW0ixiLimYdCR2rtK540thCTx
1x49h+1hFPm8oXIkUdhFwUkpOd4ttul6FhZIv5NuVrXR855vENWPXdvHQrJ2UGNQFNdq4DcUma3t
d6fKs+gVr05f1E5XPVHXc5NlkRJG5uI3Bg5tuZ5grqW0i5IMblqf5Pk9b0+yqv70H3z9+aITfIak
n9mbCLp4dkcJDGuLai+6IxcefYpRD6SjCoDhos65IAEoZ0OmNeQ9EDZxlkFphkG7FS6nFlsCe2hE
w+1ufTGjxEZZHpcqqmu5aHQ3lqoZDuetUm96dg1RdHHL0KUrRqMDuimBNHjiQcOjlEEEM4oC7pMa
5jnyXJP3XOvz/vDtCdYInBeU25XviFx5y/qwLrU6mk160/+51Q5J43Ty4TLvrLOI1QiXGuL1z7od
71mlm0+GTozCFEvnPtaXikpBHY5HY6Yubk4eukLBGVzLFo6xKZ0GBeFrk/CUJzXsKe6TOUCeqh5A
gTVKfO+IWqf8JE4FlUDJ/PeYL3/8MhPE2KouYVDZEn6BQt9CppAYcOIy5+eLQyIF1Fjy/xW0oqcM
XVtQ2oDmx43fyHGsX9XH8oiK5RXGhF0sYqaBX+5B3pstAzDLtrIvnL+GFDvlwppSOVKvTPZBlqtU
lgOTgS2+Gv4o2f17XY7vj+uAUxf9t0yACmkUDi1vd8ifIlovtbw5y+dmnErDWH9UdJ2v8av9hARJ
+MjlOYmAcbcQaXm2OwewL2PGef3RGEVeaI10WshSp4hqLZQIFax/tnvU21FUeU6VG7VlwMi7kczA
mTt8kWINm2Ktbt+bNBFeB6OoMlN0q2nqz2fMd7UOjyMnSpw6wldnixGf82h22Xa/xXJm8Sw8nJBA
EXHRLvxrXTzlvuarZbPiAfDGHmGvbQqjTWQEsdyybcoSfYKIjrQWjoOvbssqQPKKqR5eovqQsHHC
ZSADqeqgnC5XWOiSwGgD6ysP21s/tQBSgjQtPaPVA9Rrb6OmT1UvMr8Oj4qIGNp1KqES/jbzWuG9
Mp+4z2f24RDO5tv8fmuCDnNUpV9wr3thiCacvkepJJfx2VkZhedzclzeue2HFt0Mrt7MbhmtCJtr
/KcqmKQSBHAoN5wvWfX9xw9F3c78kNJ/rCy78lQ7bRHamcSMGNVdS883dnpBK6RnpTaHTZ9aJRM0
KTAJIJm4AX7PrDe9f7TL6n6vFHNtsot0cFUq4MdpuN03TTJHEx/ech3/lP/qedpIoJ0XB7tt2jzf
uetvbwxFP7we27iA+4n10hLv5wWwCSQOm7ybcydhEAcZx47myW9tjNS9ykw+SujWecZr9/lvTNNW
d1udJkFxXO6IczxdcwSlw+Hwb1osP0fF1oiRJp63/IFZAjt908/4d4lqlgfy+TItzyA9xSbCNoqN
B6XPyOkMO8eB9GSnN3WzHFs1cJSYEOKwivhC/E5L0frwIi2FRy7gbrX43k0HC1V6k//XQ2V8MeFv
hL86Zt5xn3xJ31/xjETsgL/Ya/Jwj6MMSdYQE/RGukXPNTkrB/oN4DdC5z1IxSfqeR/VO0ftIyXT
hJ4JiJi1mpCg3nGUrUISuepD3qlhqXvI13cJYheqBg26u5W0oJ+s8UlKWpbD/E2fWh7zhq/fcO20
K4tgC2Syoo76lzxFaPBhUq/wYh7cPn9UEo/+Bjakh224J/acU5r+i9jH0xwWYIFLBG6FICU2nuFD
RINXwL65Bhx/JUjdU2JC77qYMZ1Qnv3US3/3mJ63AnG23AXYXDy7D78KWIwDI/DxR0J9x6qOLQKr
H6Th8khNDOANRoT9UfR2ttF6XJ1sLRVcVapnik4nniTL+kDpdf6rpOmfGLVDA4wvDBG04+oinrS5
ul4ARMFV59pP59gSRSlTa9Pk3uCczLc8vs6OQGeAbGrieVjJoBMDKsM5nxWuxyfG6yDLvux7/vVx
ZwJVGJ5sq0esSkym9fMup3lCo+ZUeSk77RPpGphFPOZ7HbTFwTqmEk0V7bOzKE9Eq8th6C99yKH9
F0MR3V5VwFA2I73M+npnkYhkTvJS25LfcpT4tWcdbzPJXaUuBrz0I3XCrrDbwjgE3R81eWRtg5qn
y8oTvXfFZdoYkqgx+xifLFR2h+murH2Mki2h5JndufBqA8PH6jE3OgXH5NPtzh6AOHaDn8KD6wPv
st7NGP+VFcFTXgW3ovHdRlRUpX3ThiWiBwc+AD10GxsDIqIzXE8viLai3D3Uos1GKvdcnXSbGmIf
SM0g4Y3Dq4MvZas13iGOLWYdril3F6cnHrzl7T92AKNlmSPkXAvVAQSo0WWeGTbG1QWobutJslhT
PEt7aRxVVqR9olcRfD1s1/ziXyosHAizKkyYNUpzbTJN+AudrfCehgs6MaThue/8CV8GF014pVjo
GfPX2fKJVY+igY7YXKOssu9vCQZEo1yB+FviqbE8zpdnmUEpTwrKjKYokyoVTJ7RCnMCl6eqCOv+
mUNYytcJVjhMP/VWMhdnQmFIeOeDN5H7yLyNXSt29XTp3jOSX4tztrTQ/d/71fFkQ+CFHorQMKEB
9YRZPTSb3ya4giBmNom2Sf/cPeaw8nSjqm/wUmLY+q6vUPAlhIdm6nJJU3xhrUOQgvgcVDWzHIku
TEohJHKj8hMb/TwAc8g2GbNevLo/75Q9itKcV6+EL3UFqeaurSnsBRMRmyOUxdN8RvwOotTXo65v
D1LxlojWEKW8oO+idkxM5qhu/8neF0H/8Bm8ilYXeQIsI3RdugVY1rUwIP8OVMl0sryarQ/4lwwP
7tXzh8znS9bAqUVqNphxZrYkz8KwFeKZ5fUrRfKiHga0fLOKoQr5pTNmWg9M7X/Ku4VpW5IX02LZ
pMPQon82gLgV1ZXZHFTCHmeVuUnqZlLUU9IqRsZxyQovsd/p2BiGxf6H+k4VLuAhaEsdqY6j/GmB
laqRlIXDVtjvEjF00q7Wmh5/Gsxo0SCFGXfiaJ0E5e8gURxZwxy0uuFPNCjtIZQhUAE9nm6uu5vN
j/XRQpyOoEa2W/HZmjLYo75BTVH24n5Gf+gr4wBPiJ8Iu6OxAQeje/Rrt3ALjsdCT5duUyMj454p
0vrUPDAwNgAbEAzpASxVvl62Ij8uKL+tcpmDMlll1ewPOAy1CcahJahjRaf3IXEYMxhxikm2jNAc
iZmGL8KGL0wOsx7Un8vXwCCbSQmIRf2fu+5HHYX8o9riV7ktNlxEpcrCwfuNH8uQe5uuR2P9KM6t
dCdS58uqMOh1+D94zIED78k6EUWhpuBVDh3FEFK/T15nwR1dDYPRxQpeyjlipYPOXQ9dqOfoxZkp
tiPVXU67y5OhrRVTRJkszL7vOKyMbYZ2pEPhGaIEAKW5uf+L0E/JG+z9N/x3MKEwJS2Y4F2R4UzV
Iraov5INf1pzylmRbMJDWaHhTWiXGfOlW/tgTis/biw81vyMmyrInUSeEI7b/NFfvmupV0x5NP98
1qDtSKobae9mTCe5Iivq//NFJYYAnTVJt5XxpLo5V7wD4OdGznZo0BxLFQHAJ/grYcUzjOzC0HaA
0pH21coQFM1UdAzdK4/wkBLOou3jVMRAvHtkEKSTiW7z8yVZ+rvyonxl2woDJoM1nEbC0v27hDb7
f9AVQRBqosjrtwKyMwE/Y51vNFjfxEKvHWu5dZ3yv5XvbB+DTy7Za8MoBV/pvpt24qo8+LyZAkz2
L0E8yBhluJHgzw++hAt90VGbwQGKW+3ipfx4j+XB1S6OR/UdTPpUekQaKRydBXnXlN85iL2/n60m
rdj+1lYoDNUjWSOFNc/NjUEjlp4xXBCdFIfvAaZ4LFQZT2xWDTe8VZO+dRdQVosjkGJwg2m5o0Lm
6LjK6WVi3WQBDxei1aHyl9e0mb9RrwHih//P+nGkTE6vMt0yaHf0S9NZfuAPKr62AnULpsXmd15Z
ZRCF9PzJvF4NbEeI9SLkMTW8BSMrF4hSVZa6f6VkRnSFd6VyAgMABkzCbwXQ2jwz1oJcvcZ0TKpK
jmA8x5t1hSPDyuwRJcciqctAGH4SM57rXVVZbRDstDsgNQBf30uueRp09eRvHIekbTzyepix9MGd
gqTmlbszWmZO38Fh8gXjeBO0oT7Nw2BOMgpTZRtnKOPZQ2FIc0S1ThaMcGahEu5AP+dSMyI5Dda1
6jQu4rMKHctYwP5OJjGo4QSUEw1/5rOsF4BDv2rlRr7whp7pT9uNRJpTF6kmft3kIUC8y5ZE/gx6
9JdbAT3oRFILqpdMVAe1GumsWrLNXCtpXW+HhTfE4xwqFpqRulQsFeD73SASpnx33n4hkGrEpeeC
JwCsLsgVdxdtQwD7X9ZqL4avH1sVtj78jMu/JvHJzdperWxpm9VahFX2Mq+KHdR0r/6j4ghBWShk
PxQauu7JjvUjFnZDuplu6bLiUqJIqWu5VtIDBzQP67Th2qPS3iCDFt9V/UqoVZFdSl919x2iHU1p
QsCGnIJ/XI9He1vARkt4teDaemzLiTZIKYRmm2nHdUmP5E06MyKweFfYC9Iiobwp2hyVfUFE0B1b
Pb3JuQelCyJsh4ii0e3JRrmJjJ1a1y4OQ6DUCd11JWzq3fn0KHed6yMAMgdcq4UCtG56YLffa4rr
6KX7X6qb0nGQ2vLxlb7uh4hk9SBtgPxR4neLjJSiO4YIlzYLO+bme43Zd62ChxyHuA/m9sJdjUX3
dCTd5mQp8EVkkZ2E+sq/3KYg0SkQGW//GVEhNMk5NkuUpkRsHL1U4+Fmm4SXueOMhUgvnYyBf6Bm
FIb+Cwdy9qX8gEtmmxdJCWWrYj/g4qdeS6nF6B+0Cwt3ZgDIbHPnm7DfFEosL6cyoO7LxOLvFCcR
6hTQl1rzNIc4p/TQFnl2Pmg7bW98qQXQ7s+axqZjxplu4x9+Zw8zVZ8Pask09rHO7Pi28Mpzj36y
F+nrud0fWvCm0ItOR8tPhcOxA0sO8mReSZPnDbc80dcRcbHuHaN2/JCOsJqt/RLntHB0Mf/sBqsj
IEbzBnCR96cWouYrKbz7fZU5CudCzVYaI6t9kkq5E/Q5nMZLsKqg7YrJ2g3yHc2tGB+aE3N91/lx
9cPCCYjDmJ3ln5n0URuW2pOCfSWhj0hT9Ph26a1wcF4DnZzjLVotKsMWeKSpdxdmrhzNBACdL1VD
K04G7x3DxfSDprzhIoYijOThfhxCnOfI4Q3eeROy6Flr+l8aQ49/TkJxYlN4WZA5ACLp/Sr3wZtJ
X7qgzcmt0Dj5zo2VZs+wWFZUAjuOLOKRfb7S7fp7p9YkYVd9X3P7NReCsV99MSx5xC8qcFxPFv9A
v4teOzpVKab6LwVHM2o0JJiohUL6SNbfXEJLvazaKxIboLsUJlTyBpuJd/9D7dRuryjxyl74XSvD
KTVyhWywuYOAkjdJXxl7BiaCfRLb5ka0UcBt9ukw+9m+fsbPSUHx2bY2iVjko3iURwFDEEVD7tkU
46v493CwAKcWNSYrxCS3k4B+8cc+2zhVcwUta1PwpSPsmj3xOjgc3TWyA9/e7heIF1zsGpw5CeUI
ks9hYDqWUUcTUaCYYf+QLuEOZEt8oUeWj9EzBqJilTydGMuVRqkso7tnZm5r6uud9YQt5ipnWCNP
/8tppKsJreCbmoAXBYKCcNEUYwlm0LENwe94pOBJNV9q3HEQzeW/i1Cd3dErL4QxAIgvHU1+enbc
xSHOIARJ1qBgIVU+1iBRjHPYIpxSQ/GFrjtjgsmk+JeWDOURlOAs09Wdo1H37vm0VInOgFSmlEr5
duyUiabQGe22LhwrLjGh98eTUWyCNZjxgjiIi0zIfHSHPI/CPdUPWJqK5hl0s53vByvP+MFDheD9
R2HqIkWO8s3RRDfH3FaRACe8rgByiusWPDRL1LjcH5ZE7s+8pP4trmtVUYhu0tJMJZtzrOW/OD3/
49X/eMLM2inyrfUNYsPBSaNeq3Hw8IgzoyDFRnOMow4q3AzyCOVrmS9IY29Sx58oT06VTsxK0UCT
V51tNAN1BpfJ3xIarekuk6XvBsuYOWocJ+0E953E0mlKFBj65ncZZZ6jaqpK7WAGUY7XlZeOG30h
yDVZbDmi1df6XndFcjBdZz5cnNNd454b4cgbZDfA+fw3eOfer05I+2oUlDBlwSTPZjO8o4SJ6iaH
eBxaCF2E7KSXwPVePt3mSZH1giBxoLW8/E5w1UNss3QMTBwRFrDxQN/uj8IxvPpkfBadk3YMA6yr
RJLUBnQl70T5OLw5KL5m3XoNcnxas6eSSKgU0xrArrl7uLZHrWcseySZdlWbgR6pAwN20ieK47Jb
ZsqzRqdoVzMHtUcbIaiF0vBypIXn1vC+aRMnKE7oerMCapRfFYbYd/lppU68hCfvG1WltioVg3t2
HkXmsv0IjqziFWR92ZaP8ijitAVJ3nY2tGk+GUJ/d1nqzmlJBt8WrVtN0fFQ8mrpQmyTlaSGV2EK
tHOP9jgwidfWDLdDQBA8Gc5xQGKDVGRzJy06eozWDr2AMzCZDp2Dn+8ujTe9+65GcYvU9DwX0Rld
DBIQnv2TdFSLLMMFzA9RMcbWqh4WEfFgiOpEsDGKm1s5e0G8B5/pNwFjdi6JUfTg2rFGn66PFcU2
qh3OjWX7C6qBM8f8jcqqJByaDck3icERGxBQoqftJ+OZwz6myDKWt+HD5cUG2EMcUupCYAVJjOxN
ZVKziAz71FNrQhAjpwNZSPysFXyzktnPe5+KHp4uhm6xcn3DIchqkFW9UL245P9tTlJgFMFNhQ81
kVRn5vZDccE5ovGIf+nPyMLtPkXwpspMAYZR6VljasSKZ0MfQbvYARhNm3ZIG0kueFa7cvQBdLec
sYDVhJUacQjwvQlQljNdR/j3A6yq9XBI2VMde+WL36m9n8g8zVws5Adr6Aax3+DVDagmTxWOE9cg
mVaAkkYpdHdKtZJlvnpKQkQpYZFQUkt1wOijGqClHyGdC351HLNVsoU1S6MPatrSoyh5HKbybA8N
tVMuRbmm7TwB+LGhII5FK1dU8N94DBarnVSZeAzUY/W5ylUCPqDsitG+4nJgelu3/EryPVajM2mM
StZSzQ/HZr5fAc4qSQMX+jBo315Cfu9zrADhzdCrKqf/rLSdnrlCOFBOpNgyAUAaZ0u/6Nar4tiY
mKuof/bLbGiWLXInTUXM1TMK4vy+VtxwHrraGPhGUSK4YHw/7ePByYDrLxcX2X4myzknM57LMl2F
g57o8pEuGYLR1ROTTr5zbD38K7XJ8iGUJBBcIWsqYMmoeHHHAndyiCClg8cwlWKALoT3aMbCgOWF
VkfhdzDEQ77DsqF4tBitAJSWplg9Np6f9a4iixO+BKg1DWHIDMpDcUaXnpli1c5+Rn1D2bQOmAgG
LlrhLfnYK9Jn5BAt3AIqfQs/H0SPlYQufCfXmbioXpR+9aib35GCq01UQgGSljJVSEK8uEW4fpin
/w3uKnOQNevMa8s78CWbm4Uqk9b/iR9ofalnKlahoIi8ITLNpq++yUFGkXx03qSw9krMqEPS2BIJ
XWdk1KjooAlx5hXteY8rlouYRjzZjENJVn2svF7eEzyTVm2nUtngTQ4LYPFd4dU+bqnd/rbU1ymv
C+pwdzQAxZxZqCxSZNguhTPZXldUIARq+dtYc5M9YR2LZGOoYRdYT2swB78Qj9d3XxiMRRV/LR4L
xspW6jSy07YGB9LajQXXnp5gGI7mobmwh9veC3AbqpSisL7gpyK1MWebY/yhPtCQYZHO9f9d0sLt
u5ti72ahVVmZh1P2sqyCP+qd34qX7W1hTWEMj/55W1n2I2NO2OH4KiBh7i/n56fOkFC8+NcayXsj
Yqwu7AjbO7h9/lbGpgHJfct1jD847VhD1b9+6rG8cYRbgJDVOGIUwET1/24o9RFSITGYAVtIE4z8
tzQfNox/aDQ18g7hqrCL9nHYmhmTwMpFUYyPrMjcCBCoXRBmSN0DNqOmZoSKHlPH3E7dtu8tjhWJ
aFf0SP2YeA9bzflvf1lx3sBrhRXEK0nROIHQDQnZoFuNp0ixU2UxjIbFnpHOCozH7FNApgh8tBj7
Ptw2FbgeUt21r/mqCe4dXGJ2mDXOPak2UgJrZCGI/PAOt0Nigx4nNX+AINM5PyDwyPXOfGlYSH5p
OV0xktMW3v9imEi6IUrmUor2yBr6cbfrqQHnpMAGB3LfM3X9p8BxsXnbg3a/IBkD2QKBDh7/rbXJ
5FZuIOdKSmAhZuWixwzP3QlHmOY73HJRFnE+RjxkMTSH2lGQNY1Ry20cdhAP2MAd9yICUwF96Q8f
aEROFKvWL6OFmoixkpccbFxKonu+l/tLpUCESHlnWwXrt1Cp9O2v9Fe1Ll2AMBuuu/bLYJrvJzzU
CiY9Ccff37dpnlaVB7q+GMKoNmggTVtrxhuKH7ucmHVAcw/PXgekcU7ogRoAIw0HwxivobKIhzek
esVNs0uAYmhxuu+5d67c1eAAk6Gy2PJmlolFZmwxouTC/zIw3iNd/zDvHEMtz9urfOnslAaYM/Q6
SpAbcQse02LeZnMf7719FYE9GIg/6Wtbz2KqLpzAItGgBghZyJP/ROurEzFcrZfiZ61tYMEoTr3h
VHpdZqwCvc63I53Uv0m/4wJ1QtLIkehq+UhmKkeVpR3SN1IU96/rYAzZ/9nceWCwepoTazu64+mq
h2fTE9qIDR5KNHWuwqUoalPiIcAo6M6VMppxmYgn7N6ilouyuEf3b+WA8m4hXn6tjFP2ixHYvJ21
LH/BNjZYg7xF1Pj3YYIW/cYLaFvZDBBw6oY3Wxn0jje/HwF99JfZdH7qfAH8znQ8xTii6hZkhrU/
3/+0xRqpi6nhLDqX+2aqLREtk67aiTglTiI8AdyHrNkpBpmybk+8vqvz0b+ggtz3HHm5jq/FkeZy
P12ZlKZ7v/9gXeCSPsTL/vsubzkKwzKCZnG90P8DWEKEdTWYFDTVmD81030AoVzbsQ0QGArtfp2U
7oot9aEjfI0JXVoeEtObMbqR/86HxWJGvdszK5RuesNDx9vlIzQ5qu/Z/c3UxVaZo2QfH4zaB1F0
t7f1D7pq1PQ3eWOY/kDpxZ9Frt2mTrpHB8nIFEiXylv/Ixp7c3Yk8UUQ5AyWUNxNLvnwfZs/RLLx
RyezjXAaIpDKNuHOSjPlg1Yd8jOsflA3Yx7nKgeof24Qq9+9XsrzU6e4UtzSntuUVxFwHS1phPAs
d5Rty0oJmDnAHUSDPKYOjgGxcXid4sxSmZDBVQle7hox+eurkdCvWeRs1IREC8BvbsGqLJtXgMof
XnvarqDoisl6kIDtx39gGtKNPtdoN2ciKXWod63VCnJDXLyE+jlfCg7gsbfwW1ZsdgybH7d0E5fx
GVzDyybRe3/TAuBDLPG+eeQkl5hqci53Zo3/6Atv2HMuN0xv3khmCtUYZrlMN0rwaXK6JwouGlB0
BcMJNT7mTaMSLw+ilnlnm9QKFWl2NkhsoNNWg36OVmewAA0jA77uFSpfwYcD/goALOH9vAXB/n1/
+0yWJBebM2en4/f82/MVzhDemcFGLZzWu+uLuQ2msVJX2uH5Nb5j704NX65p+jmoWtLEvnEYQu/Z
YuIUY3Lc+UzdvpMjIM0Rp7jeCD8++VUnrDvGGG+zm27lcC1afddvsAz3KrcT86Cs9I8vPmZslooV
oJUYEAdhtXmZDRDthss9eD/wunzYy+qfRcbqzdj0Wrp9E0y4izZyaf+vXmTQJ0wnk2aBsK8CA+RO
ziqQTb0WK6VNx97sJmHZIShI7YwP9YnU9ZBeKkf1XXGTecyGBaCfRRzQy3pkUAiC5YXvFiCWLE1I
Br/llOIxa+SY5jvLaTSR15fQagKPLm7nlkQZv9NFNDAuOoSJQ2/GKAqjfrTOA2cEc35kC1iYsO+0
VLdxke2LT2o83jkQbvj4KOSd5JPGByHW4qtPg5BHkZIwCKmUtauBnZujX627NvQ+uq+FSAHmRL/k
vE453R5bOIOjYbQqQlZJTGiFBuskvCL8vlYpuSKc1sQNCclC/9vfcGi5S9dxaiqQgE9nRAdGMMNQ
bIZWMz7G9TWI875/oDtMAwyftUoaYXVPIdc+prj8URUja0xewBi/dAz718zmR0oOrxazAdJDqGYv
UUcEQpuXYb3YNbbqSo6wyNyzPL+hRKZo3TN4U19sLzxHMUOltv1C4gi6cahTSWsJRTO7iSWrDJGT
o59FREUmfoQHAa5a/SEJqeFztbLaMcqMfrHXITKOzJYGjk/H16lLheCivasEceSxBOdW6aI/Kq9j
ZdMKuITK0NWRuWz0rGxHkXFcD3ikbhI0Cn5vlGyzoBgQiQLkAWfIa2pIsb5KnX2BZrQXPAbk7XWI
YK1sjhjvzMmsif7Zq3M5BFRos3Axysy89aPkGraJNTDy8Knr2E2ZKCFzX19mjSMCxVGWckFTvKkk
lrz8NrSYEYtcjTwrCYJcXToPy2zvJMDDbcKuwUT/N9eZbuTbb9hswb6iNE0UHopqLJPuPkBLxb+7
avsajRdCnr4/T6pUx4UR8jEX4nSAaxrhd3L1nrf3C+4POc+euEhv7nbRlhplj7EUZu9qgrXPWmad
4XHFwkP1hxtBgY6qg03v+1TY1Mj5rqRR8Oq0Vh2ghYSUlBg2SN9HAENAMwntXdanOuRQuItiY5cb
j/XAyRLk+QjzzpePhcyk6RifPnaGDWKGByPtsdzdgVAzDqFbix3ptbbV3J7fMPhECrf8srROLpsL
rKpGG3J39iVvZFnYYFV/aEdpl5oFSwKjvUsP8Pu1xsX/DCkB6NxaYoEKuvASyQz/TtcB4INPBTXT
9ZlKQskbiTZB9/BSHPPffdlPj2Bkr9BpDQTkRQg/tn32i0PgZFGTNRYN5U9LnRezAz6wsZmWbtUy
FsdFh2Ikl/VCMQwuv+3RcBsJgie5Dcs0j+owAjQ3S0S+LVhtaj6pTsG4Vg/1yPx2NgcvFW92h9hN
/wYVPZ/SRaDqIe/Pi6FVc0Y8GZsp2RcP9BTy8fuOe26q/5qYNanXiVkVLiBu2vdsR7w1l7oGSp4O
L5QqBTEn44XdWfxn2cLuKpjgvBtC79r6usiIG6ufc+xOwKifK6eu68Z6kGqo3Y5Tnj4B503Uhq0w
TbBvgWEXnSN4tLxLB/n9qoUz4VEKIrwUSIv4HCxBH2xkjblSiekaoOhLgn0BWdx7KegiyBWBoEHV
WyCj1BJy9jFrCfTClWUsO1JoSbM2D5dMGvTiH27aTUIUNXhtpCoWrRHPgJOWCrViqpZfmM674yCu
YfKIinAfdiEurDwzn7mMM7ndgZHQfmX7XMA2GVd+oAn+li6lKb53GUyNNrtPjFYjC7gQOddALg75
Qp63fFfM53XdGMYOT03bcDtOxOg1SzCFpsmsr5ytRR24Kb2AUWw2CGoOu1C5AhTaZYOcReZ475du
Cd1DLxX2asLc3GGLSjn/aMkYXsqXbBMLbqwFD7iENF42XsUzeEQNnYIJPlNn5iG9zegHQVz13RTi
GacXFNEr9s2RJ7UU8qaRv0JjjTN7UghKhlaQ+gsiOQJye9yr7KhBp9StgKDq1/t2UoMJgeIjupHp
UORcULifGIZt/F4IMW2xObEySgKwkKDS7bH6bJjiWeyIRrWc4FtIvsdCFD5CbyaIM9Xb23akJpVc
hXK1hQyxWaVlxItaKelpDzmByy99INUOQ/LzNitXt6mZ52QXjHJcO3IRXJEQYrVwDBfm8OoRt17i
B0r1DBBjfxor9wXfKGgvzHWCXEYmkFAO7fzCEBKd4NlSQhZl+zkwtjRxOi7TAoCKrRCWnMpyQCbD
78w4QipyafHWdAK6VVgvS/AyQi/ddyyhgNneeTc/p4DKeoNrmf8zUgmzAPGl1lFZ7f8oIOQkHEq8
Elssc5YwPV7R8uxQLTwHoAfaGgZSHrbSrEbEe7aMS85aKHinQqLPUkjvwIJvHhy3Gaz7Zp4wgMUF
hqLG1NNnG9ATA9aEhkk1RjukrHJVxn3+QHW/guZGkbKz/0+Vs52P1BJd28wTCuSmheSZR6zf6CUN
m1c2BvZuCNGCLrpAMd0E8fAHALnJTBmfdABvXKqZsx3zvq9IoRrUlBE/mc3Qe8cqoWPL0KfODsmp
imf7sX2HWtV7oTd0La8PpSKlo5zRTOBYJ3J8+Hy48iuPEcpM31dQjeQMOyMPMNNYP3BU56HszKhj
MUCYgCBVgmo4mJaO2A4U3CpU2h/3SGrjSnFnHt/LTReGx8j2a8eCPP9i6RC0jGJlb4WhIqhiRdPU
MFoRSkumQ385t5FJiVqmkrsMZmNVtV0eRtsoaEPjCWHbKPf5mASgQ3IJ1Qxv9ZbhMROSQT1N6mA8
UyolkB2TNqyoEJZdPFKgFK8wonAGRYf9CskEGVMkLg6zHY645OhGxt4AyCRZ8IBADA43+iwfQZIW
sWist/JT2H9WTpSNLbNUWod15ln5RiK6fW30kKUJaZwXpmRJxqkwjpV2F4jWDppYxCm9Lzno0JcF
ipLJjjQHiYrsQ7Y0Cx6Wqfy/uXs2lXIpZnXV+ZedCOJHJBTPLXlbBAUYIN//nUJQvSCBerThhTLP
6CI+pOC8zOHfObkyMNnnKnojbB5ryrLV91la1TSeMmzJs8HNtWpcdv4LksOgzupjP1kTpyXFe4QD
4yXBSOABD1SFShFgkb19Tumknn8PDhn50/qEIric/m2ZrTmn/ZaglfpCDZU57rnMAr/aeNaAHz/a
ccfNvqiBnW7wWsSWmEmGbab3UQyTdDzwKcpKLXq/w9kVL9UPpEX3b1d7IcdR21NkmTNNW4EZVutd
Iac0dTfKGXNUKEj6BuVdr3zAUgrDjSjOhNxjNOOH54Viaz+3OnPLTvCpmshwaG3s0G3XD3uM/TvU
9I6vVxBd6EMvsfl4wFpynrfUzGBMRI4v+gQsFzd4rH/jUpm33fjDjO2WEGKIUapa2fIoyVkyCFVr
/yLYW2HT9tYJw5R/6Bq0rMhEmi6awpNrjFxjq80EsHLRw1QHTsaFCS43EG6BfS/8sgN6vSoZrL6l
M62AmRBjKulCn/PogXI8vb1aOQkplj2LzTtX1emM84rBr2/BUaBR1gzIpahHjaM9XhPQmHDjzL0h
pvPPJ+GwzS3VrRVNih68FQXBexrG76jiNjgE141pX2YL29AEFPwkQoq0jkh6TSSFWLwnKqD3UUuP
YIXZ6F0xlBzV0sVMhpp5Qfuv98gFG8RNpr0MMMe6SVehDvh4ooWqNxyPANwlmqQKN2KFq+kwiDS6
R+mYIpsLpXIK+1KemlGx77Yn1HnmgU0MYxWawL+nWuxuj8PzK2c5PciUlKTum3ZCrZnzyMVHRoLB
Dqq3W1BaI2hlhF9r4+WclUq/yQttT1485RBhoakjnBpqKMV1ZVu//37VZQxQTb/EtQN8XgF8IrRx
OU0RPsbVjyIfuJaXMYgFJdwWCjQn28ES35J6wjjLNTbtysCyg+EDyhksoteJS+mK3he1ff+5+NNz
GO+HhEpZkLSu1WgyOFedhpJq48n1L7Xf+aJoKsCRxzsOBURVh7uWoll86blq7R6hdbFNfwHuDD7I
YvdkRZqXbYFHQ3D0idCRGaEV/z8Fz4ZAjqTD0iTmRKdvOjlTc7hK/eNOAu7WuXcsN3qcAfpOLO/e
XeLC7Yo5XvPNeQVWNFEAjsAd0G1XDpdTccM07AIqxds/q8r21u+K9CpOFBK7bldxLmYdUT+RUS1h
bduvConwMEbjaQ9IIm/cTQXoDTeADcJj2Urc/sLpj/sZ3rQfL165aBZ42w8OhC6Js7y3eXYndjh8
vmR+oZABIi59F08dDDxgWtlFZHGkJwctOi6VZQ4/rfrSfghOp1UTqkLGqiB+BmquRNdr7o6HiZ2s
XmzdDL4KXik7FmWbG2H6X5A9RzjT4F/QLvYUXbKbRIAkbMnSqD95qEB23LAKLexdXxyqwuwXYxDU
Zijqb8wXgZpVUsGWus4vUB0ICwgIrRo6We4B2mSNOoI2WbR0r73K4rTAcf6WBg89Ma3gvmCyUqK9
ToUShkcWpm8obU1kBLOoKGkYKSqiRZ8GWac1fsAD8JZwDwr2VYn4EqG1hsGCzvobpm0xOqZY1Bva
9/CIxvZ6vf7YJtZJ0tkhk1OZfCx0pmza2hi2FoQcHB6bhaGXmItXuznEDLDBuTDtbOIr0EuQTJfG
wKrnrpWCw2RTcEhzYQiZJ+H5651EvHht6vdKHJXpSEd6rlSD/2WYEve3gmbRsyQd9/jY8iT+S6kQ
84HHKFh9H7eUobAQ6WcWPOGLP3CnMmfnMqv/LUruwnpkhSvY7YpmnckvJ1Y/URIhe69ZyFUftjSL
lEaHRIuUYHqW0JC4+zBwV1WR7/cJvCREnaNOs0mqLzLutRLKt1v5o/StgkauBwLWhRNjNLYZUn/z
xhuJp3Bts7NWww/BROF1TzTR5ZqUZ7yCsfXNaXp+pBtZIuvMdAWZAZxsyzwo3OK247EoZqiwAbjV
+kBPET49FeQ7TNI5wWLHKcuUr8do08yDughtA8wdxAtGeFhwb8qAzTehdJqYcs0skhwJqMNq+xPJ
Io1U+96CFmVA0tZRVa/xhyFHP6krxh+3ZmPByAIJ3tbjhjJqnc+jHS+QCt5JjiCaLH6TmHTFogho
tFIjMvIXh4frQCy5MTcp1VdDhR6mqXJ6hn6q/eQ8pPWoYmNCZ2ozZKwa7V70ZSXmHsQjtiYPlM/D
BQ3x+lH3uDLcVtDild3iDDzx1nlCseSpCr9JRp7kO9p93nkPk+57NDZc3Z/SLTURmeYcgtD+rDYG
DoW1uJNxOL83gqwv9H07UsWSnOaIGQliFvIkc02k9VG/vz6rEFMxHn2P3PvA17j7W5Z/RydObhBi
Vug23NmU0ilSPILUwted83rOSww2WQmOAXiIj3DwmIvVnV0aQM6mFrlWYpx+htFH0KEvwXsYCkOG
nK84HOwMU5+8x75YkRhJiMoZv9ChpWz93BIxANi2J8kqOi9jLO61Cd2PNoJqNsHPhub7tSmNb6LZ
eEV+lVtoL7GdVJiREXoqkHT7CKrZfUU12WVWTQQqzO1m8bvEx2duT9XUeuYCY0G2LSL/qfvDsXM3
JeF7nKb0mtVQb8++SPrcbQpjyoIZWi4WTVwwZpcBg/A1AyAJN0gUR+Nezc51Qh688/9I/WyqqLMO
VC861dkYdUTJ1UNl3oaOX8DgMoyYUAH3XkFW3YwDGt/mcDLbrAxtIFJVoeUmYhi7bzDZz0q/gdr7
PFmPHd674+rpEKBg4LwAXW4IlinZLc1JwFqZx9+toLyaokkdPGDRsWZb027KbVLbx77SxpmTueOw
asiF4cjowfSWRzVv8IqX3jqNImBB4xgPm9nBiUF77ymfNmk35cyzrvnVYTQpGtvpyWkf5TCpZU17
LAcczbGs2PVgpJrnoUyebR8d5GOOgFEX+ouCJAVUlp4J2SFCFCgtKEXl83pe1L+R0HgnAVLw0zaS
8458Of7oAPErSTg8X6yIfn9eFzH/G5ZkyrsG80bUphcATBtZcKKmNUOVeHXnOTF970MHwvhwKzjh
OmFs8zNVYIAtC/rI/k9LekObONHf+7jzDqFplqqOTKyJ1blpgvGbYJGmzArdmlG04pq4qGu5uuxk
/sZvjhXMM8q0fJLOoYK/GNmKwctZyaVqZ20lj+KRgTixUCchFQOkCADSOJO94tRdlIVekSTrDEG+
4iOnSTHZU7iJg6hfP6Izr/Ua/CVEqp78KA5854PNijN3vypdWQClJnRPpHsLUsKhLVzCWCfje2pD
6WY0YYoCNaUVGPV+GrZOhkxmSfI3xcqdW72BCgBQlLn5oDtrEn1A0fEYgYVP/PdyICAuGo65eoIp
idbTcLoNasLB2EgUVk8mQLIOsZ+OAX6ht6rUBsSAaPHE2v0CU8tVxjPP3coRupkps0lhA8cMfVGX
iKFBkW8zVPp2qqxA1fA17io3hjN/T61kAnR6BZSJhZeZmAIbfl5Mr+ns0RFvkGNtQfm7xuLlpIOu
NjGlhKhL7dN7IvVS/TqissV8tH/qeSmwTUKf+s3lWSKOmSlRXJebjJVQw4M2m4+Wkeqvp6sJfHfJ
oaPUZkpckzBiVJ8Jn+OCp7b3ysNFemPSqTIIT0b5nkd5ExVQx3o38O0QdI/6FSCEgAAJKWngRWKE
T/ZnUZ6rs6sLgTxyz/1W3SgFj8maEsztiSbbEVlz3b7Bz18NL9I0UQ+3POptymOnpMTiAckodtEo
X5mn5lHpkKoWV2wJLZGf2mUQZTBtNnf2DHht1d0wUgESyDOGyx2zzEqeCyuQTjoIT+3qDqwIzqI+
mSP+2H2rlEULAbHwPBuI/9tsElNudWN7f43UX44MnVmnsb1Jji880ZA7RF61wgsLQcXeyghZw7le
f6tgyMliHMOPMIjMR/4fjLewiBjkppXi0O5qckQG+oqyJbbS/wCzu3WnCLb2ZZUf+TM8k5CgiXOi
ic/smfF8tvc8tLVelf6cBsOdVPoE2Yei8e3OUJhpmm0HhURiBEOtqrYuk8Utxy5fb8ki6/RmhnF6
ZEe3ijss2atciOp/PFc61MUBQEHLs5p77OS0w3BFrLDiWUtkrBXNMgE5zxVrXDlgTyZrNoLpWDbv
VoI3i/8IgWY4dnPG7cvQGlsDn1AoeE+mhY+d66/uOCGpVrT93UjNkUcoPZEKeJQYYOA5APxbeYD9
4LVHDYhyO7Tp6PuHwP/bge/TCfPxLSxbirwOYdMnGRuhKDh72KxFP75FHdNwq//MRxuVp/JhzKHw
nIWphxbVUrXoI/L05CsKjOobk0wdjQTwJ7IL5yFaVAHgaHhsxq0lgfBJM1Yyu5XpfFM/Q5+q9DSi
iamwN/jo68mtRBNPPueKFYoD7iPTDV6Q6TCyOapuN7omdYcVrcITCZyqQBOzEek5gD3EE/ZAGdul
Y+AlOjxJ1L5S7j+yjPVkiJYpmJG7wR8frcJ3cKNxJQGsFGZ9JZJNav+Woi3mKPFvhsrxflEfTgrt
BBIC2c9UMDLkEwCcUKYinfBnfNJpYyUBp8jqVTwPEWkHEjzDPIjIG1PSMdIsgHtxDKX6ZawZ/9oI
AS080q6MZsXSg226KAfkapDW8IQFbGys5smu5q26A25yGm9io+XxdtRXpiQ3sZjF6RdSwSSy81ya
IVR9XmFAybikfIw5xK/NKL/S+2iCGxWk3Gk8di8MMVaK1Z7UAifgZIJB6ubr4PGwc4qcDVqrOWkz
FyqD2TiXHfaxaw4T+tPKA563FEUBancUqDFimJRToHnOwDePOiQ1zfQaiFij0E6vb4Js0PuwENZK
PhjlfMqKpJlBnpupTV1KIInsjdFXQsj0TEEZvRZtY+Dxh0KyCVwBzwxqcYCy2Y6QVv6yc96+9PbY
hnNisGCuY1xyfAXbT6UprnMDOJQ+He1RtZb/Ebd2aMlK+PK8vMnt0+hbEwvBYivZZezgLMy46nHS
9QRptu0U/qPDBxo2Ox9VNunGl8Qt1/VKWUpt/hTuE/n3oPGcnnHdYws3UcmO+G/GZb3Z0A1VcZN+
bKd5aSyj+B3njucRlitsdcXIb2Q/Md7Kld9Pu6cMOatverQ2DXeAQfx3JiHQutCfUVqtgJ4dKW2O
SuB+W7RyGuMUXWIZ2OFiHNCmXmuWWLm178vwEoUuRh2jAz3bKHXg6YSC2euyHRwupVRpEcJOeDIL
/eEq8LihTwTyg1gCgMXUv7peB5f63XK8klgYqQgJEzkEE15CbjnmbpAoEX1bM3ORpfGyxTrI1EuT
n2M34W6bpfWREdrv6NbQipvk75k3WVuzgrywGGBZsj38+yrkfhuHGxmsCU/JFGGQzMHMmjOv/nEz
ZoMNO98b7AO7wSETntlm2aIb5zY9tXskSQ00pJXl7l0TWRRB4Vm17z+RxwPWMbqU8CjYWg5T3ZT0
2eaMqca0QI44nLzMNiN1OSgXkqK/gMsNNHqgjRAViE45cTd/Z9H3YHWZUMvkHiv5bVUCBJcSvzkh
3KclJs7fqT3OQrUmF0Cw2JDGvOcM/T1AC4gavAvXdA9p8E0A4cErdP/jMSdTqHHT/Jz8l3gDY1+5
w7M9QwE3T2rI05czBC5fzKngJSakpwB9GenZvGKkwqjAWfhboYSHwA6IuL6xg4WAM8fjikBBoNgK
TicU4qKCMZ3isg3Xw/ba+no6T9ckDk0o9eeNUXqVNRtXytkt8xxVCwyWKtvPQ0RF13IrZNn0nEh8
qvn3JrYO/Q0V2GWIoGS/vgPFexBevE6+wKKYXyJTuFSNQvPrXMmTC5N1J+gu9YdANdWEzCMfBL+I
x/j1FxILWDILvtXWz5aDDWENO6RzZj1NRcw6HjrS67J1t4PcaLshceT2oAebiuNOIf62ja/wmn7O
39bLwTe/htC9+JtfSV/NI7/EntsWpBlx1FLnTqNZrNDfQryVWOBkca8pd3bD9wxXnQQq/YlZ7rYa
kzC9srGO0aqUElxhz5EO2vTd6ZuLCeVpk7s97uEJ/RnWql1X/IC4HkYD1Cm1VYFHXp+D4UYhIwTP
vSeijRNeuGee4qPRtApxsGge9b3JFG0Qxr4/EKGEPakPt+TY8WNeDqSMGtd6geFy2vasweAcH9Ni
tmu2Cxf3ctC4ovKPyR4ZJXh15cgt+27WpOS4q2MfppwoNjm7AvH/TCdPBr0PDSAfXcXDjzv+VK7u
PNLVhiiJFZambPXXdrZCzh0CjuEsJm4RsRAgm9S0SOLlScLpXwvylr6qBFl3R8SuW2Sx0VXJ/KNn
WxHt3GjcRPYUBEl8katBVFDrPWppHAss1UYIBGl2LeYKqCeILdqRxAbha9cw9kQ0rN6PqXHugbwe
u0m9ixQD8QvtmgIn2rJ/YKlZA1KVpMk9iby6W53rekGqnMUbftUkOYjxkpaVpv6lL2lCHjEcSfLG
X6Lg0YqdeeKK5yshjGpddwdxK6bmTIJhGRupxNLVPAHLFhlHY668TFyyR4SG8QfTOr6diqEgoRzt
n+VYkO1jDta68Fve6U6nSdPqoT/VitCE57cE/+mtpcqiezR8io9dsZhlOWdxsSgMWrbtz7GajyrN
0TkxcMC6MLozoyycKYCbko09VFyOCvDlj+Ta+7LoBkAPYbtsWQ8QSOIinlgWjLl1f240Uw974PWe
aB2+TASI4bxxJht9gRbxOIAnVnsLGDYWzz65UAQC7x3ynSjGhCXz3DHpIUKzTIUj5QFGlqA6epyP
uUAFb4V32YZK1vWQ8ZXL2GmRd0gVUkXqxVZfPW99MqaYkPRHYuoOjCdqhZFT/xTgnEMKNpBqEUIr
FpuET9A7qAHmf3fZh16zr0jJu7Oy7SKfsJvMq5sKJqKkloczjijFLRdKXZK9TT8v9TRM8H1noENz
AzYq+WtudTjQZ4UA1CLFJsWw09tzS/JOFNK5UlsdrIXWaC+gSuFEB/fHs0ucoqo68gnE5rcH/3Oj
qyynVv4+ar1gdZcylFgz17DUgOpyERJcDIJYFpaSxtg0HaZ6zSp5Oje99okUdcvPQSZZ/an8ut7D
0UWED1y9A5Bw7FwtgOLIMi8Zd6j4UfHxFjubSHDbli5X2DDxkSnm08YpQee/SY1R1xm5iBhyiD+n
9PRrOrk5JBGqke4711p7L+WmFHRUAWCuOxzD5Ag9Sccgfx6WOBOUXEKRlzBQaSwzPcuU8CfF3ahB
ZudNwU1DptlbFv8C2x5CO3oZfG1dxK2hJ42lmSxZFJVGVgOgzzQR3m7Kwd3YJDac+C0uj66w8E7y
itK9/UBy/kl3IL8JpDDVm83PI+eRmxQMK8EkGD9+b4r8jNXql0frYZgimPUMENGrjAJ8xTMhjlfj
mCS3Fcfsvsr+twSF92CXeL1RKWv4t8TTsVchBljg4Qx/EnaaVWDDxX3KiB5Omdu8RPcFrfT5LPy6
DzMbZI7sWCEu+9V+/r4L+RSaNCoRzXsagXMqTAWTVAQ6Ywgi6BR0n21zan73bDTiR4L1JD6v+AwM
mzzMoqd/KoOfVg0SGcc9FfxhmHc9IDigSnXG1lI8vusfVxZuE8NnKp+t4p0gQIGdHHaHoe5msE6Z
WwVlKjBNTYgSZHS/rBvwcSlu6C9o0tyZ0wYZIanBUNZ3VBbuUiZmHZf9QoFlgfjno46FGnTucENw
jxRuxLnfc3A5V3SXUwGRxVf5FWvLuzARNlvoAilbhqie7eYJ+Nxfhu6ZrPZC50xZHuHWPP3XRYxx
oZ24yOARAn/crHFcY5AK4Hrwwl9AENY0zQyqJo00HoBLs7MEHnmPac304zi/7lWlTZvxvwtm4+ZW
VBqiNF91YZZre3EaXT1dUuFKMnbfDQxp4o9S+5s6BajHZ4wgWifXpuIAvzT8rR52w2AfTU9BaFUG
y+2FDGpG1+O/u9bmRAbxyHcWcK6/H0uB+SUCMeJBGtzfxKhy5WYBnCndfqc0PAe0d8mqOXO9EIYn
NvQEaKumNwlx3ajpPNQbxfNzRsxnQI3NIa46H+Akcz4HYKsEn58Xzstpuj8yZJIwlWgVIFY+6/1Z
hjZ452aac6XRIUGrIhMru+6hRsVhiRsbr6ZYo/f7+c4WMQmw1lYgho6iilEcaZZzw/QwhaQUnVjR
9Hozio5s/DqhDJFBTsruEGGtmvJwTU8EPMbgaOsL6F8tDJQHQzySXLoLU5xePeqCydjVFvWrWhWn
lxxX6E+C9goAF0O0w/CxiZGAgcqdJRhx4wI9JIH10IihOFMAhxiiMLsJ5PQkC6PN0DmbDIlYmGce
qMhKzDPr5Tko10scJrHxupjWSUNeJub8ra1sHrBbeKs92Fj8Nu793hRasYgoDZ/bLBe1C4bjdNN8
kKIYCvDQzL6S4LPcG5q3Bgjqt7bh9Qv+i20mOxwPwHmzaoOVkd51XUmNpsia4X8oH/RQL9+f8ZFH
1h6VmuxyzSOjL1+7Xqw5X2EeatKfXBZabCQvx2vlmv9+S0XsrmE4TFA+vaVESWF9TEYSNWwizltL
9nPqBvBRC8LkQHxGzUjYxTPazAV/bquu9WArLbvcCVZQWd63tF35U87nMmn0AD1F/K7DDmAgxW9I
BRCDzHi7WJb0cuXLknK5tsgtfhvJQLOqbUoBGIMhqpSaWzIscca9+3c9l13OZOrWBYdu0RZRhlvk
oPHRtnP7FtsEkGnDpyrsE2seHnqJg2XVOCa6Vxh+APnndTtl0YtIY82du9JtM8SbJkT7ow5xF0lq
Ad6/apUsmOLxOI8VAnZZwG2vGt1XSmE/IKKzR7wmuJ2b17yKiVNdzuLd5kTLfa57OznTW7WvjQKY
4b+it8CyCusni29mNwhnsENJipR7BXz1EgCVzc+h26SPfjq/aabhJwNzK9f9wQJ+TgoqqXH+R3Ic
0YUpdyiWDW7ONuVbmLJu58xbo2CeDdltaFz5ngKLkRdfwRWkcr7yw8idykMzDN2UeNNcW9GSxhEH
6P3+MyC/SZjgPh1KdVLKqNwrj6i9Q/EeQpm+RWxK91UsQC9/16P/WPDlGwEqdWHiDsZXl0pjewgw
PfX1L2tSBE2jOuZoeDB5Iv9t+UbDXZVL+DbegYnkUheidLYUDcP7KbbVtH8Vmc0nSprBXFpavNTj
STooF2+X3eiFfZ9aixPT7o3dMsE0rIzuOERucPE8KMCrYEXmyUMawaDtOUkJ/tksg2AKDJlyWW8T
E6Aw1nxXsglGdkEgMOUcJZi7I/P/kiWm2ay9V3pvMXZS2yrirzMU/YzsSUg42I0A006eLlL+YP9S
mLpGoSJDqgUQ1hc7tr8KGt5BRHKhUbBdZ0qrmAfatR2Lbuy6gunWrXQ6bFWQAlm0zTKPfsAaIE+X
mzFHACmqknCjPz/wklQ7nWJOa/khJmKQrsfWRti/SDtLFmx5EGM/ZttfdG4gPKam4P4M8UsbYWOQ
i6IFYCMFOPAgfYi9cGmyOcx2DLAl+2yy76tyz9pzUTJzsjWk9kOgsT8BWYRLem50uU46xZDabwh3
gUoVWvY141Sjmrj4XUpxJCVXALQmncAJ26fMh52o3yaYy9U0kUQYwTMjUA1cL04H4EduNy7VLSQL
HAinoIinkr3fzLu4J9KEs70L5yaCUXEbb/az/216s3oYUEyIAo6C/z36A3H7Askp/LN60hGeXklJ
GkUfGLK/mLYulzOd+8w2MtdNeq72Av77ZP/GvmHUO8UkaLgg63jDwVlxTYotWBUCpdDf1JVrmhDv
l3H7B+vX3ZP/82tPkOz6qOqSn+c4q8myvNhamGVEYf2HX7Vk4F+X3ahZB/DpGS499o2b0MeZgY19
t3D0iZ3T5WwbEN2ZpzRBLeUVtB94CKXw09zd4qyMkBZn3ZmORcI98b+xG2wwLKux8Sf0kiFX9NVR
HDay535NUx4Tc4wGAmba+3XeFuJ0jwFPL1ggMwVCdpkbC3D8Q5zmcnybH6+j2bWoqxTzTd2FVmBF
OpGY0blVwk1GD0BSi7tz4mYB4liP+8WTQ2Xa539PhV7DRb5JqqFcH2r73axd3JB+5/MQBLS46rTS
a9jC6pdkeJyGf13P6EW1N6MM7QBmjpi77OGnEW41XB1VymUz9Ep64opuOIXLl8ODcMRjZKEHo8+r
MynxaDaOee5zWi9IHM4oiToZJ15cqf+nmRpfVcrAdU7S1jy2oH0VNfSwXiOEAdN+nkBAUYcV7364
sBGKL+hLfMlKnybfzPC54ZLbRFSo9yf5plj/YH+3nXNxuIgj0JDHCRw7OEH8NAsSEkB6D8GGTB8H
f7a/RS7pv98fWBIdDLE5PiHv31xsll7AIIXUI9IBQJsNWsi7G69mmUWFO4hCtjYiIFNUAfBTPD9b
pNx8T5TkUQxKtBiB1tQRwrAd36Kyu8Q7UIBOV5grCoRS/qj1zd/jG3XuoCEa2xWfocb2GzAmsd4m
BwbBO661V50EQL0xHiXfZZlRoEIj1fbc1tjcbvq5tk9icHJX6G3slov3sKRY4w7T6Oqsopf/ZUFS
3ExUI8CMvS15T/zlmT/rUWU3lI/Oe16oCvSdTho74PBOBhVwlCTZFY2G91XjACBg8bZC2iWgZRpy
qWV1PyTJqvTyWzOCPon7vZkrTl6Q6VtcCT8Es2VXMXxq+jjdTKKYgvFhfsF359JrKgE+bqVVM5gs
8rflcRhmiX9GILKwkePc0fxXOTChN2/ReEfoszVdnBWlgoMn4Q2JQ2sCKn5PezrmEBBbhWcQvt9C
1IRjDynSR5S1ys2VE65vL9DcP1oMo55TgIHVe3ArhytxAltRO2CKZLj244nKluwPJrPAs1k3RmLt
zA7deICTBZPS1mBaPP2vM/PK1JCVrL/vZfD3UnTRiaLmFFuuZ4Hfr6TOlOGpDRAkA/qa0Usv7IDT
2jZnNZ9Urjri2UMYSWcVybVNSmX1Oiu1cZ6+CeJdeTqOMg0FHfuHC2FpOK73v1nMOLCyFNsJ/Cgq
KqrKj9KOJEqLoFPlr5w+zndaOMOqOOAsp3QUJNgAKKYmCAr4Syd17CO7dH3KOo/evlQf6mbOvAVI
pmkdefcSKg4E+C8E72wbhM+YWk5No/1wl6j4//UvOon5pQVnGlEUhF0VmwirYxxeap9KpX5xickj
GVcYPeZ0HEk0YfY69FROxB/afDrpbzgwNLDaNh72SgP4gpSGzRSrkpw78uVHkiYQ7YP2PP7SbHM0
f5lrk8X/5saoPD2xNW51Gh3dTnJWy+5pMmvzoXALh79tpvTkntbK8jyLke//QqxJgBdU01yFh1Qc
/LH/O7A1XcCeujn6KlxepHlMXP+jXmN4upbxSnCW9+5WsM7oiQMp/Ad2HOd5D4m517mJoVNpdXdu
o5N9WWCHgx3A4ZDXui9/qLP7/ReN9ngFYXLowaFGGtpUPjgv6q490u6imS+nA9svOdoyJCFl4rZ6
SrKjTBdoBE9snq8VgvcRim3myDe4fJeYq+H5okObyPZqrtpPpOYBv2KMUROrrG0I1O+NEqOTf1Vd
z8ANbU1VbkO//jfs3P3gLur3Dle8vMuR6r+q9TQrEu7BOQe1OMcUsL0MEcz8qg3K/fYza50ZIRU4
eVBigVUkqaPE18jd8u67QmcpEHsmTFvy7tXm16rLx62xMaxSeilzXE+6UjRcr0ejf/QJ986hgqI7
Ve7L2uw+Rqgqvh9q/uecwQY8UX4dEOf/zZbG8ivM9jv+fG1Bv82bLrO11l0lFacwJbbsZBEWaadz
6bYOlIlXA9IwA8dbqkq+Bwu81O9V8XnEsu5fkh7FPJD8juGttxY3ylBKBo3umSnh3GgLfFUHj+wd
Sno6p4SHVjm4zcwIsJLj5d1OXOUOoSPzU3x6CNGDTwjtJlJHcaZLFEG0EewUcgwlMwtj9ix/MuVm
KQuMCxw6+x7QiRFRrarH3XzAl7duIJ5ZvPCyjojqhVDTVPDLApbFNwnLBtwz7oJhBafzgtjI1Qc1
6y8XgRncZIrH3YD+wON01HXD26Neps/RvwmMVoJqpEH/JuuIXQTBN8bL05ddmEZ/ArHG6GusrgqL
n9SSSfGfE7e8u5nEXcn++Y/yxceCdkyS+VI0idJEcDtev80aaoUr+Bd4lkyA3iIZkggcZ9y9epXW
Z4KHdYF6h9HTUZrmXil8aSS7e68TbbewvI4D8jyOLpWN6JE95DIIK2ozEfLYOa2I2AxQ+X4tgpgE
VBZdmqL8NrBRGtlTUOIMIh0a3DYl3FM6PWTL2REKfdyVhjuGW/WXvmT2TGL3NY62hhtuGvYTgdQr
r1wd5eV8yl4KIHp8sntn58RojKcsIdVnvK5wAZkFs26MtDPUfrK8ivsh7O7ejIxuvhqsP6L7HuWm
HFqhQQhFHhb4OsCWkQBruSBV/IoO9LPe1tEf+isOmAaoiRgLktV+TugwuEChX8o2CGj5OwWxqwPm
Y3iKjHLPVoKfO36EFLPnA7qMQTClZzpck+m4A5YojDfNkkmndA020tuUFNIjuI3NFzcJPJFL6YUj
KO+RA1MbvQmSw98U8lVD8SvgUTQJgdN9v2tjWBkeBV/ZKpxGYfI+Gg0BXl+enSkNg9OOlUGcvHj/
UA6PxjNSq8hAxlDCzDxKEOwEOuNGf3YNSch3MsKINcCZIgEf+nEbkRz3q8DayzEQuxYFcadZ21ap
QnIY1T6BB+81do49YN/H7/g7BTMmLd1gfMGZM24X/FE1E2DHLIk2oA7M8JccREdwnXw4OjlToMLy
x4Mr+mB0tUndPWqoeCoiy6lUaXdx/ZG7P5eGcTOz47pasmqUZtDGSu+zdA+u6tf79QwZsdjkDQ2j
ThvxXJxDNtJDsjo9jmg2N7XaT/B6BKK9hf7G9hL9XcYlpydy1aVLXNihlBCQMBvN+qLZ1jT/1Ve0
ok4PCOioYF6hjnQ2zEnjjWo6ErwCgQP28uZQn7I4u27PSAlIqzBjIHJ9Mubwf2/BdCVlRhd+3hxb
Ju04LDreSM2En5Z1QgkCZjfS5Jc/jBd3RTvhfDCGnYb0UTLU5CJJlyXppgq/GrAcfoq6wt9OXrrn
t3VJ9cdefihj6O5iRSmSC3g90ukNefJbXtacVppaCy4f9JDbbil1jqSEVO3o41f+Mgnm2gSsWMP7
PJISxZAj5VlR1GgvU4NQioW15Hn8yGzDbBld5y14H8HZc+vVuF4nZYBWMAB4S6755Km3TZZNAVJ+
R5ecGfjJr51FhyzwIzyGLVRidGYykc2QPDJsZiHf5UYhJfWqjjxphGa36RBmoSwkfQ6HbQMX6FCK
qif6xF/Z4hISi5izhy9BTIFK1m2RKdm831u34W6xRdu7amLx+n+eWJxhPehXj+hOARB1US4XSRQq
V5mi6xqK19TAXECqGXbzbmbwyHO3YhUVoSHDUVdous+Rj7GpozIMZ8wT/T6GKFK1iTuWkCC5NCa/
+uH5D+wKV0//iIb3T9fEIsuD2V8S9f/GSEi7qFMrJt6rXmrvdfEEExXm0bQg654isyCzwvWDU4tR
5hWv/00deuffLuHQDDj1Ch6BIvW9o8/QZWk8TPkNvIiDSv40hdfVwOdftVDu8Kdlf7AYe0Lt7tAK
OLMdxAGbwktodEX3++d6hfh8pOzvlIexD9RFU1zPUVXJ8T+4nxhVdlEZSQNmH4aHxFrU28BBTsaM
g6MXZ7JArBDlVXntwTFBaKXn5prXPnCBx9VwQZyVgmgoT4Xa9DB/PEUdXoBlFcCvj8h/vVc0MXhr
qV+Ig97IfkAmFFrA0Gocsqdfh/BuKK0GTuLoaZzI5MTO6RJChIAGe8y2nafzZkWXd5ppQrMYwW0W
V6EKgCM4zM35c9op0EzNEfAaWQFkSKGGoEkfphEnIln3aaBm+Ef9Qk/pKVO8EH7ezzVWcYI1htY+
/TSEVI7+ETgbCTV6nZ15QGlfoCYzrjuDcw+kGf+3YANB+a52F4WQtIgUvMX30H+SZnzbjGhMu8mI
jGnb6TYqQ1buH5DLqpWeAVWqWi5xTG8K1loYG0kkB5hURAIJ+MqmxOU5Pp7PEEmor+v169cnv+YH
QcFBDovCWO3ALmNI13hOqna/0PYtwx+s1mDkgc74l8xULDzRjhmgJ2sriWanSrrk0Sof6i8wa7OK
GblP2IrFKMZrKWhXoEduDNHswE1q7AuEZD9063Sr+s5d6RjOCQcxXgXe6rYGSYxZVRLFU/Vy9VET
E2N/sYdm5NeudvTMA4Uhm3LQvfTFhxwLjKxN4Cf6wrr5otc2PIAVXPqjeVMYa0WVTznpLWolXnRp
QpY5V0e8l9dEAl1ZcMk3LXtYyZDffBWYJZNwfnyiZLiHqwSEqalDwML9PZoCNAAOL0MdAUFEMdQy
NDHmXAsefFZdJAm2V3J490L0/6KZTJ/OkNmYgs8WmKzE6tQSL7UA+HTWAofKgICJFgnlSFG35i9O
tVscrjB8mnz6dEo6PKl/YzjFHMGonkYEuNCtMouWlOWI6onKP4phrAp32ntLNe06xssHZV+Q49iS
8pi/vHD0vX7blBJIymfM2krOjluoSsCSrB766/paaZ1m0Lm9pr/MHeBqJ6L6/yGgmAPGm4A0DbDt
5bZcL3tFZbZJXPa9NFXpwg4oMnMjjNg60oJ5fNKomw5l3MFKon5qP6LGV7QutN3Qu6uUP5tU1upn
kYsu1HuD7moeTneq3FWCzYh4Kmu+uLlTIG7ov25xmkUObLfKODq0F2Fz4lDjzxZpqNBVZd5WrQH6
gWc+CKsJAsl++rS4woI+wcRwst4dhtS+Q0Q87t0KSmUJvAN7BQdj5WnBRtHx/iFEYdG493bUPsZi
3HVOy7qHzYL2v6SxRnP6lk0tDsZOTIij0QejDGvSzZACnhmJQ3p99RiU5M+lXYZSwtpKbsZFC1h/
ls9mVAhSk5bb7ipm6j+OmY/ynh+oHH2XzdHa/ZytinVNx2HOjTS4cd555UEpOyhMWaruzMWfvpP+
TQ7iiEU2EShoHJlxPVP+q7owmErrCqv60njX6xtY+E+MiLhjk/j1BorPVUWfqs7bYmnmZHrEmbrL
+BYMM5T9Wgo1imMZzD31PqDuZNfGqfOxhYShEyO19ef7iR+JimP++/sHbwZ8K5MzGqH8zNzgq74U
LPDXbNv2R35USaFsbD/wZM2bRSmOwJ3qiLQuvmB0oYhlIg7GvDuX6RGAVz+Pw9zQuKXXiGIwYjZd
6OjkEezhcJjsaDbssjr7LznmhWN510xPRwfHOZBOyFIe9rRgCuhABFTH3wZxAgyuc0Y0IBHi2d6m
jZWsSJu1yCTSyQate8YHaCVmEq7BJwdZN+1IO9N/Ta3YkPQgLa9tR29sWb0wQKtbHu8hmIdl1nuu
LRhO4ar67Cz91U+hKx2YQObUhJaA9bTGS/373Wj4iHVEtjwVx/Z9aMrDMg9g5m/nUvSELPw/v+zR
rwlNXwMCeKcfojFqdKO7yX+fcJQx0JRhkpbDt9fbv0iT3SrYbb8sBh6xL5kHtSlCepu4RPpwCG5S
MLb8pdG3SdZ+n760GRRjVzGruaiMjYVlc082w4VcTNyjwD7dxZgkzE9a95aRxGLWSZdEIrM15soe
v88zceo/jhtm5hDmIFEhkjIl3v2TNnCrQ2tGtwXTFKSFQkWp1SUlS+zSl1rYo0XKyXY88pyyEGFo
mDNsoJkn7CSc6hf+Rc8SE0h/u9h4k7epdYU/26D6DeNvyrdR/NgYTe96jrZWgi6i17NcDMmvFEdB
oPLiCzSSa77XjthN3JZ5XhOGaKA1VHrJNG4wFDDoQxHWQztiY5gfUsskZadkLr/ZS4RiCf33daK/
vULhu/ZOCPv/NBSeQgM5ZKJkfQRmB8cfYCi/hbuMEngvp861MuAvQ1zcYqC6CxMRGF12/IlKJM6O
yTgvwwFKYFp3V0cU/aTcCgm9JsF/eRNosOreFQhwKqh6j9P3ru/M3EIkMj7SXqgP/yiFZaQsQPV8
RDR8FHMCEXxN2P8GMLz+Wyxk12521Hwrx5BNLGndjrIW1ZTewBZCFJvgpiTnH75M+GE8tOpOuDuU
4qyVy6Xb+Fld3sheal1aJB20w+0TRL3Vyc6yYY1x7nLxxm9P4pIlfPSY4uOog37zBaN9gvFohQQt
qutXvvpXoqSQEfc7HtKNBQH9KMuyBoMf9EbeMXX2K012oLoJzksyul0sz7fIre3XsFhi4DxNMAP8
aiEHumxZQOvESwWMwTLjTpkKWiE3PKrlZL3UpCeupNF81medv8qppZmt1QrgchQBnaa2znYsGcXi
6FJR9KMEgIItQwKJdNM8w4yaL4R3p8oLzxlbUvB3eNphYpG3VkSFCqKZQlrmqjWJF/NYiRQguPzP
k1reT08EOl5REfC9ruUBROOd3BNkhnkrQjahliQ1nPin5+MwrsY+ICgcuQ27ihtIBuPw7d21Fbtu
pyqQv/R2Un+yS3NUC/u+/k4QBzXruueaGaywc7hMpQiewSClDXzHUau/hoa9rS1mstxiZphhXxk9
cJtIGG2abrl/KV9u1/hbbg6a/+I6287FapxPaB0Z/0CY41xirQ2s5PKjCy9xUkBLf9N1oANZCFgw
VAWwYgRT/oqucMdn2QajnjrvDphlNXD0EazvwIHN3y5fcQRuJHC+StGbUN1Tdt1p7ZR8kSAcaRxk
B2Sk2Pa72Bc88Yp4/U/PZMhetYGFrgXgwwfkT8srRkCfJ8luekQrq53C6SJWjAW21G6KO5EInb3u
62RGY0zVoEUc7EqG8xENK/wQNvkJOQEG1DWZq1LVpRNBTDrURdmTCIT6wJsOZd3kgS2Pw0rshlIb
Rh3iPcPW+Thvf+9JycjCefg0cnV/GzXEeBXPJMi4bPCkd3m9uQeLvf9Sm+vjlrsUjtdX481+MxPx
sT7fl6wYmlTk3VqyCB2CvDRQQ7q+c+HCi9Ylg6TkfTOQMtYriFYCNZz8K0+9yP3q6dbfgu0pLBLp
ecmaeZFADmQIZfsdZOellJxMdO5SzBEy9AkOYvTthfzXsQmD2XzYdu7+ZqsNLXtlpgKfJc8M78XJ
Cx6s+N6Kc+quPP7GxAKjrgnzYJqhQ480xcB76OUBBYwyGu8jwn092X+x8eH+IsHEq10G40DW3iHy
0hAJ+Rm/mLxkNXhdqCnUBu5R8CsTpLcZrq7hLCl6rKe+L2t3lmrKhtF2yIfNkrjdfkUfTGrMQPvd
BcloBsC6OmmKShzoHsOWKQsx3oldKaxHLPIyqL3VTV/3e7hsdgdZiew4u7QUJfmLJgc2xTzO5KKo
UCR//cNlPS3SyuHOXTS019+7GRlhZiHlqfnsOGOE7SeUUaLCjeWC5D0Lq6gikWTuvUhLtvUqK291
l336/Q3pz6bfVqjpLTvIXtPEzmxqiTrEt1r9RPTm9yZn343zmNFx4oHX0fjzZXJeGrnqucGZG/7h
gqD2ijbhbXcBXnD1sWG9BCp1B6iJ5Hw64+AngXSpa6wb5Z1fEbXvO41cicR00szqWZ8sevC+ZBaQ
aONlzbcMrhWLAG4EKQx4fFQkxqlWeIexFR75EncZ5qgFDvGLRgePfZQjFnOOO19ViduO/Sha7mEG
8eQoWAGJP2qvQasIvXSw2LMPQ2qRa0/ElBUcFc2Zl1bx3CVxOiImR3CGV7yMbJiaXxUZ/lPoRvEt
jbjXui/03eFWS8JQ+KcS2sIqtPnF3gbiglt5zrazAzI7EWSaD1BqQdcnt/vyOi0wFkNjHYjh0oJ6
A1A65YMZgemyAf41GHpFwTQhUY2JHvGqnyyxnHlLYsdogc9prScNG6ALlvs8CznrB57uV5IAVgmg
9SmOsc/qe0kYKyJuS1Xpy60GKPaUr1Yf/in27CoI2YzhgVXpjM9sOiV2Z46oezc0euTKacf9gnyy
VCoePRvwyrm3GFe1/7cvcAXrin1WmdtUNqcEQUqJSBnGtUynihehynMcxEHgKAoGtvd4DgdfcPPj
YwX8OSioXj/4vqvzISvjHrBXV/B4Q+jiplGaRyYgfHILM5MX7d3ussbmdqKEFxdB+gCJgZhoAUiG
AZOMhnsXpNwTcdJDOnIngs3IBSHSHzzNHOGQaeC/5sEOeUKsakChbGkoOTmga2luAFxXjm0qQSUu
CQSabSYBcUli6Lo7O+3ToousOwhUD66g1UscwLFy4G9gTluwcDea56o2AZlMuWfsHKcjFSKKR4kv
S3c6MzrSLNhBTdkmSenXgo8xVbkMvWZ7gcqe8mvv1QnfWCCDG3qL5iGGFltTK+G7/VNn74MGcwT9
7Md0goUyknq8UhE01lXQoNW2Jg9awrbaEE1vLwlJq/xKY4zizDDi8MhMVgGFOZUY0ZUoDQEa48Dv
H31KiXJVM6IKF8atAk0gF+s/scnUuTZPLumzqIDH9uqzjcQUkDuaNmF3+rzMcWe1vDBb9z5If4tj
QNS3VinsGnH/h9vSxDPZQe/RvmNh+eVhMVj/kF/VCptZuedkFlxx1i9EBAUWCGFGbdr9mbcS4xpx
druzgKEZceT0/TG8EoNPBilKOlWN5NwhDogD0eJc1XGPurgnMpGaNZmK++33fMBH+JcbA9Borz6Q
aSW79izGgiKVJgh7JLfmFPBKc3w8cRMgPzUa0oOCd//VcMq7HirlmMmknzfSaXYCebJtEQR7ex18
zpqKYVpf0ZNGqyD3a4prPniPghuAuQu49s/Vi2m1Ye48wHaRQP4/eeSL4kgQgOz4ss3Ti7LJybHG
xA5Val0VOTGtKUMTpDfk2BBF2W1ZsUYlvoYV+843Ad/YZZOY8IeNONP/+ffqWKeJQJ5sliIjt4pY
JPq6hAqcPk0CbAh9xeCpZLDuLqCecHL7YCYfEy73O9N/2wD9UScTEBLqad7H8arSotDml32O+bLM
IhS4RYy49XwtFPsgFDqC+n6RGtvnExiOg1G6gRvgSPTRV8NsDlE/Vg04uF5ysaCwGGiwKhAxkVmY
qWx2/HrFDOzXiMrDamDM7joQ5f7d5PLtu0nIHtMPj8hqxH2dv1VkYJesPVIalKAaFrb6AHxo4wL1
t6cwKuX4QBCRMg4o9nwPHwGYrimLkoitiyD7nSlJQhiN6wmZFEaFnFZ49MQAlv+n0F78TAFYX8PE
KqX03/9HSaYM/lM3uILgoAyLQpKIZFzLWeWPTshrqFRX6G7rA1GtFQi0wWoXGYYj2Te2OT97JeLW
m2Bl9avNL7tngXz4qwS2ilBa7FpD38ESeaeaW8rzXlidqtgvGgzhTmiWEJmtMKtBxpr5H0wePoRZ
hAwZsZmo2nYy+P1VOeZM7n3RA24zlaS5MTzPH7Im+Uac9WgYGYpR7kzkFSob5eca5mF8E59ishLv
JNHPI/qh6GOy2G+Bqu+6RMluTiKu7QDqbU1zHb56IjX6uIq7LqCIZ+qXj/zzNKGY9LGZ4LoVpSia
tSDPgyraKMk04kdaxSVaTW++PURDLG98L2R+JUUqV+++g0dHQKd4fQ+I/XKDkyeaVIwWHgWoPgvw
uTauMBkoUn3h4PePWN+/oln4luCvVmyxpQXI0hzLpWbWpHcnYTecr45tZHsow1WeMXGf3L6lorJh
Ret1p4G05O+fsRuRUPXNSk4RuuPKJRzGun38dJ+sBcBykdppcg/mQFVmPb7+7XIHcM4h0OnC34bU
XcucKl2IbuSfnhCtQ3shtMIrXwJnxSs0UNobmF2sh7zshbRyxz8hWtIoFK32lykUeoSioiRVG36a
cmdduKxkkYqLG74blZ6/9fXp05b0l7zrP2yQBY3uht3uj0kN61QGl6I47f8nK+pCfAmeBOMwrD1t
G3FBx6C8RcMCHVU4rWVpu0F23Skd+8dnmZQIBGsgpt4PkU7nMIvzi0ws2QdAyc/Ny4AFDqsBfN02
V0TCsheDJVluBjfaBW4G5OJWop/o2WKFlI35oXzQ0EIvzI8NcUfncOlh8VJRCqkpNopSlLKsLP/5
52iYxeAztiuSj9KWn0uni8DuohnsKlvXc5IXXB2A2zdrhTcsIX86Tfzt14O2o+oxENzdSOU/v8mg
BtTWqpwp8gjm7zjrTfZhVL6cE7oMWKs6zvBu9WqgN3c72lfDuUrJW/IcgkXCBHqIE5QcBuinw0aH
I+ZrI9PUQ9HHe5Fdg++Ig9GjzCF0c5toTqUzwmaTtm+Z1IFDtrx8VJoOmH1lgwNVGcMSd8MVQg7C
pNft8xHf0ehdYddZWibDyuPMVyzeVRkh4/16GA9S8luToS+OzgIS1QfDiEiUVo6+V2+TjFzB+Biq
zsKdrPeUhyWertdgj92ZhbrVvuZHbpvanffeYRssG4pl4YF5691nY3XN9E1lfTkGu6ChQcMz5/WG
opjXnhRcQc1baP1AqOZbW5nTJCbmHfifvtK8CgkR1J3uQBAK7SxSH8TGoQTUimehls/LPmlxwZ+f
CKE2P52rIQo+OCvfswV4K1OSdMmbm4VxgV2Sp6TyYymfJzHigU8PnW4oIFSOeFYA0w5cH5oSt9zO
BRC6xctQBe1dzCd181ypBnneEFaJcB6wXejRwwcXtWFbirgqzd7qkb5rnpR9FPvHzYbvkMyBt3fG
EIvuemYRnp+8xYNS38sB26eolb+WC0mAewyf4WPeAEMrdmByRBlRu/eDMpkQYVKbTMN8YsrlRzrj
OVGD+m4fH+6vLNMDp5rZHzYL+jZKd/AnrNaxk7MbCGbZCLPAo9F+fskcAq/MkxfagTdXr6dNAQ6z
V9U50OmwmCB1UJbURGrVpeYuoogT1ScQu7jvVdD7B6civZWXxwSpCK3+eDFIyGDN/0wpqju3nZZH
r6M6T5NvZrbeohjpheTCLq3gWJ6JEkrZEb1xvx8sTF+CnE5hXF6WETpw7Vamc6dudAZIKaiRUpPX
IHYKrrp8JjD/oWuOKRXltCwZj9kdtQeMx9LngDb75Gh0RP7gO5DyAtT7X0oSg0QlYYon6gP9dZL7
hEvwttTqFahT4xb/kkc3sFmfA/AAMauq0gyVjbJIeSNbTsy/e5bMTa0+iyD8/9sPK67sS0Z4p4I3
eWedG7r2UIj5qxWHWD0id7J8khV5noPGdoRYs4kJRPO55O7NdJHGYhn1HuoYy4fA4VrV7jHGR0i6
Mt9kJioyePZcRtASkXprCehk9oyPUtCUu8fUAlbcxrjoRL50/Ia0QSZ6FQyCQAV+Ktnh1ncMeMXQ
mDfzT84smNvzEgO5jflc+i9CjBrZbQI91wjoO1MM/7/qCgtKwTzNNGYkl+iKKYCxxwVluTNGWaLi
1wl3Zs9HebJ8WPAsZRo0i0HXlaivmg97sxhJs5sz9FlnOq09Y6mcsSPKpak5m+NgyEgZZvdva1er
zzIsoP0s0FB8Q4/UeovR7i0+rEAbWUJFHsIyaQxZiDPS0B0waF122CeV7r5hvdnjmbHGP67e/cuF
8+i+IT0zO3tcsaApO+RQCLYNPhNXpG90/Dqpl9/FM+CdVhkFTERgCfa9WcTuVSe8EBgALRaTlJ+B
ERQt+tJy9+6beYTzwF5wS/vSAlNrCqso8wpsDfvYRLkkVCB0KxO1Rqnz3siZQVozj/pZE9ml45I8
b7d793HJFqiFTQHk8R5AJDpXdmZvgUPqk4NYjtQ72fmSRZGpEITXr1NLZJ1LuPYukeWxGfBUpgm7
fRBL2AGLKj3OkrUfE64qzKk0EK4kjbYamE2U7PYjlqUxAVMihZen311ZlvHk+seYpm5lsftCNu61
kJC74pqQD4seq2qizTmYaQj5zKRqcTahJzd19cAaMSk6zHBXrkji3eodqphaaCQSdgCFzWgAEUgR
+P/MuNeT8G8jrhkcL2p+0TjUXy7plsuFgvedLqmCywr7ExNrxQDR730LiqHDHm2qxWL+HkfLnAu7
OsJq2hFbqBZSzWvX3s7/F2r7X2Q5XeJXHt5qblcUvAMM2WZ+sF8S2i3BuhC949Z3wcGVtfzXsCl3
u9ry1qu9Ix66GA8oomReKZhb+attTh2CDq0xxr77w+3Xg/R0ffvHPkx/zmu/12eBcpx0++AG3xP3
Xaysd30o2UUuj51Y5l4Ic4WBlpbzpZOPvDABAC8x9mDlkLdgCIhyPe/P4D2UHa7EAsQP0/4T655o
YvH7L91URHZgmqhFH/xDRlGxQemzJpjiSbTdUNSIejmz8HRVAJ4gJgpNiv6QTiCk5NGA9+J8QOlo
1U1tsN6sE1vCIkyWjdUTUKo1C2apQWRIUXrCbM6tIhORtX/9o3qY/POONHamkSnY06fz4hIvYy9w
2RyDuoMmgMWfOz5qwz6ybdmzUhmVNC0IWiIUagAuzq2+Bor5OxL+CPU6aemmj/B9gV4VIT/xQA4t
wbtCgRhHrgDRMQx14Z49844TgCBQfbW4s7TS/2idhY5B+smdpWD54wlc4SvgNc7JaTQmYsJZwXOb
b/MQsh0nt0Tqnqs18Qk/j9XpCaFzrTBXSDIsGqzD2HaRjrkAsk4HomA55oZ6P3S4t6q7a81dyYKV
1ytVJ1vp1A1AZY3lYDL1yEGQSf8Ol5jit4jyd6EVxjqazE2s9ccNwc5coOs28PvVej4kj8T1DqA1
EEvwPVoKdSFFHLxqIU6x9d+DNli+/OqarUqg5GnPkWbxlL7mIUkRCYxZnscAw8t4l+cjmOiazzjI
xiIN+LefJkMtv7WGHUx4W+0qvhd+UXa7FQKzeFcNJX1znajpqJ/dB6w3NIczlaLZEZ37WIZn2X2S
y0r2/BU68QA2oVbdQ5mQiYoY7cWVYfAOUnzTMqucd+9EE9gXg5y+Efg9eNAHIfRjvPn2mtVCgU5x
IW7ggjiV1Qy4nP3igWkWpcoTi4bb2bpL2FM+5xD4mgqDALBd3my/5t7RHSC8ntULHltM3JAWSmjn
iqeTzW4fC6R7hWjePjHX0Hr6YKPxGN/PY5daC0hzDrLbPTpuRM1AawYZ0Mq7A4SR46mEHW6ymjjp
cfUdR7sfwjS7gsbXcA1z+2IgV3ki/F/6LxG8YzsQOX+e4xtMRlzEdqjtgEGxee68C831K/+O4K8K
RuuKOpknKNJfpKgBSLWWuLwy2dLP7Zyxtf8amaMh8nh7+bgut+EOmZ4e4OspOBHPjtB3Jd0l21ul
l1bmPpQo6m+TodfE0lRweEO4RQ9x9Ilpbx8QrlIx2V3EzQSa2pBdAiUtWGbT4MPwnBspLpy9QLfA
dBV4jxOsL5OJUtDXg+ppyAKdbJ/Jr3mIQNmHhaJ3v3SWoOv+ZwRwM1dgcSK4rSmOZan0SmRlMj8t
RTi6BGstOeFCn3rPqRtuDQ8MBRzblly0ydSJDn1skW1PPeVzFTHchTAXdgLQx9bUjjCGixdlnQ1n
VJugqjvmhhosOntTzhVRkZlCt/Ek9x1tXWoGQX8zIiYfl4PfzSCt+0H65qF2ncU/Pik4+w/cd8K5
gCyHRC1L8LOghCLZpQBnE+uSAlNnJKNMaFBhzbr4aTVJI3BSnVFFKXUJTyUsqgueEVJUUlmp/kn4
TdOAU0gTFEb3fsMarygM77i2hpYXiI0DkZqqLdEa0gXIkavhL9avAkIf8yVjxHbNgBRSKX/cSUb3
cT+dlqhKwSm7LRtKxNTrperprtbsEQxUqzp8e+LmqLlp4WtLWZpIFaJl64FqhDIdrpScU2csbfnI
ClZeT59yR1y6f5bO97kKxIuDINL+xecGfZs30hPuIm5taemfLFivh/ZFZMYaSq3ihPY+l8dbw3NO
JYXt+4HsEFDweWFqTxSC76oKYVBNc9RX08aKc4kzGOLT86bX0gW9vixL/y/H0AooC+mtUubiu25K
LnLSd1jgiBghZ09DARYbUeS+rDWUDGwvgYUmdCliu6xQJqfjwsb03jGtSrxjmzPIRgU0gncBjU5Z
3DmCeRpewpk2a0JlfThpvBqxtCCjC5McqAktEswM16G+GdcjvwGBiCkbaXtvUUzuGiMl0k8o+XyF
rpW6EZOK6QprcgWC8dCYjkUcK9NnGfdL/Ob7agEGoRBArtAIWHgVvlM0VSA1Qf+TXhm1AnVEnJQP
eBFnAacDWqjdTjjhbFDqz8GZyCR2bfaj1nlhj4SRwuo9l3VyJeHVSM0ScXffF9sht+f/bT0j5pLB
CRrN3HqDTqFg1v/Ba5oomN8G6xTtOhzwaSXTUVV6FJyzMn9h6y9l66qYSy8HklWnlfD3Gnd5evUr
91mrCiPT5UvPf4tuBUGZIENZ5Z4xtueDnvSqEaeDEBoV8GOnUSWDRfpM7vrhdfY2vAY2r0BSR8ru
11Sk/p96cH/OByOL9wualH79YxRm3eo12SPwG/Zlv2BqeCOWjbd3qqS0j+6PZ9qZbrbCHxi4gsze
MzInVJXc1FtcLelY7HBOoqcDyKdj1nLXjWDBk2r9qrW+DxhnJo0JYgtjQmhqKQwJy0h2cQ/kQqpO
dQGGMEjZTsb7SUjY8sqyQx0b9V7BBDU65ZJa2E6J4BAodyIeXMLQlSxCx2BeHNFvObaOG4AdrGCG
jSXK7m1qLL9k/L7VbTads5hcsZlXGmZ/VD9GqLucE0/5h443SqnVPV1hgahI/YYs78QBP7S22oEb
9+22XxYmT6VUcJeLxUASnBPizxBMcwwqXxMmEWIc/TXT0bfYocDIj0n1umQRQ0679DMf8NLNURhQ
yXgAk76j/hyuAWzK3Jn4u5HmeuTUDXIZRBOiwqLNWeSxKPfw0CaJoNzvc34Khr/bSaGbbbmXwCO9
txT2kfKEw3nSJK6rJXWIMU2FmSltCAv/9C1wZ2yy4+fCUzk9RgRaO4uMzZlVXxdKgJq4bnos1HjU
etR+y6Gd6sf5Du4T4ETIKzevVID90ur58Ce5EIB3xqz9nZ8ZvDdYWtxASseVQNukRhUx9eg/bJIn
VAnFzd/YYOPaKOGOd4gMO0IbtGhADatdVrFLYn3inGzFiQ61fUsC6qr3u0Jdl7ES43tstZvNmwgc
a6yXlqG8VqmCvWKUn+7ACmUN/PLGJFrneiaKkFJs5pkMWgvQTMiQg/CfcDEJxm4ijTCLPeZnfr32
WAm0zM5WSJEUZmJTFSVJRf1uIABQAkah0GGdmUeFjfXd2t2BNHvHBp35rw6uGap4KL4SZf0UNyhW
Fm7CI591C18nFJ46ZZ/3Utl8thlmCug5EPMEX+UymASM3bcJKB8U4nZoHdjN6SOuryHA8D4Ava7v
iX5J5I2iYxlXbJY5mkcs8XyB6oFoWYhWM9eHfHaYqeFMvC7TgtUYjY0Qbt7VfKfyzTEovvZq2//E
J7eXWZMrNgU5VztHFdxgJ7t29OHvHQVuNLZTAE9gWkmG9W7ilTfK2xJBQ0qRa5DzGsBJAOAvxoxA
s4lmYGb6h9rgH/0KbFQWOfWxtfwnM04kt6A0zLwF55RAqIuZzCeVMRvcJQf64gTm3xbXQNIfGB4a
F4eFaP8TVj/SVVti/AM/4IEtbG9uf5DR4KtK34pMRmtaa2cAM/vw0OKPXfdjHLqV1WifQG8aRlch
3Qi1blRCysgcMRFpew8CM1n/EZjv38Y9iuq3ahMUd25DcvRmQSyFvdemit6YQfpNChdFHLq/MKyx
qFeIEY7z6+RHuvOS1AcnU9x8/vUC/H8yhemQ08oZgjjXUr5XLNm6Z9c2R/b9U3ndFkjnxcYMqMzu
msBdgteJATJ3k/cS1jG06IWscsPsj2GKh64tJHYJRwnigf4kORcX22dnSN13+QtintV8lb0Cw68s
bR/CaW9WgqXAGEWLIWdyY4V/e+FbBoyHjyOEMbjY4CHEj7cD/ra0T2kMX6CImwzUgIuHftVpuSx8
nOpqC7KnzpYoIE02rX3ktJ+2NEv2eOkRELRYYk5K8W96wcSho+UCrXcEl0uwHnLhpuiirkl/BuWz
LgE8uNw8kVvL84kOqbOsDiS/ZWZYLNMKlz7nfoweXtlCAzwZtPy1djrUxGpCDqtvXX3nTbGaRB2Q
JwfPq8EhilRe164dkctqdKrxSiRNVQbmd3vWwtSP//vX3OlSJ+01FyMAAwk9w3FY1dc5Qg9d/h2T
/dG9SlIIuWw4eTOYIhB4sZQOVL98ckgnKn8PbkvafcbqrcBKoQtlBFdpyIeO+VtwLzansTvz2k2r
jUB/9Jg4PCVscHIaCeh/792dsGZ9MEr6A2pc0vqUb7EuzQ84ufoK64FoYPmr9v3O1ZiE68EJLSLB
bRhPUNv5v5QObdgp55PKwZ75OcAENunfhpxnNme51o5r5CDLJF/LDpZAHihpn0jI41Olcz+6fWhi
yWTLO8uylPJF4qMrIe4q1qxp+f51dPjJXiuLVikfx4mP9xH3XQlSnxZ8qcGWHPhYpxSQRd+b2q14
MZuiZNZ+F/eR7Pd0ttaPUSZOocJk7RKGMGPKbe5xbssS+lGKvXTOvIiW+LDGF905V+40cHgWETpp
bYlZ7WKKluRDxKZvPFK8ruXNY9heuQHyYCe3v8oYpHlAYqskIToc3lIlXI0yUQyxW33FdjrWiDVk
OnsOzLzVCxbl8DItuBwPHjt6FE50DabIztqZqStO6S2IuCYUwNbpL0UyVejjK7WJqtU3XAkg0rr+
ekgBeaWI4bhQQuq+Q5nKB0MwRlai3jqCTwaCOoL4eamQH4jURMPgZ6aGpYjxUv0hHRCQwXThZpXm
FfLkruyB4AIrZsNe+Ld2mcxvY6QA4DgHqRpA+lgHlRNNLw5Y2idYIJu5VN0p5PbUvEtphlNIPlDX
th63ozLZaTGXVBNzRhEXU1ygVqTVHOZdZ2ofnkW5EHnuxwgJ9baHB5z8q/zC+/FmHE/AT/GYRpyL
m/+mVsABqN/z9Eoc9dqfS61tlJjpqj5S3MxKm4om+x1j/xCGfqWMYDV9GJ4VoJ/Om66+LKtqs4Q6
ud+h01tXfKe1lAXIlTh5+sX1OzdOHDeeVhhihUsKHvFhFoMRiJ9BBetDCaA+VdqkTQGj3NFuNBZE
bINMfbAaStVU8NQQ2+PfhX5GyBiGXyA6D5QtS8SjAxREkNqnQwOfNQwaADcpX1g0Wqs2Ik72wfV4
hHn2RI4GMzLuAcxTTxgwqJWCWbZ363n4jM+cVhZ39SaioGKTkU/EV5y11E2jI02q5S6tFqBNjK3r
yFjRqp/qu4eBPBXzx6EB4nZ+KqXnIsiUtpyOSqxIilMvQQFggRFbkef+UcdrDo29MqEoudiNJl6p
/Z38a+bqnvq/YmYw65kBmOp7F4EkGyXUDjzdA4wXvo/JHBEqfxlkTD+NZVpmRjaHGF/9c9ctL2yi
4LQTkye7kDHx43A1kK3xpEP5S35qUB2fG5JZdK5C53eLDicTNuoJUz5zy3l+4JIAW7JhxtirRgem
e9aumThdRmpR0kfDNBTPkOusNXNsthpM+8bmUCIN3Q0uF+S2AxltVUQ+fhXfAXBOExr2WmixBjEr
Tm7LzJI/VWMlIXsEIIdt+xg4LpaF0ddwqfnnRnF58obfuVyOXD6IBD2gUtAovStffOR+v/wqh/6q
NOEFHqhqlaDIBJ6jcMjhp5Np6HzMon6CGzRXZlasf2Tngzv3TimsjL8CdEkZYhoT8tFr30wCTjt+
NeXiMoIXtduh3FrIutG/C2hOGOLfi9Wlx4cMahNMd82ezOKT4YF5phgQNVBuKPj+3vKlYkbJuZ27
ginYlLjFhnFROl2ypY6Zfx0a1Pu392B1gO9EqFnTJvE6R6KD4cZB3Ro0v+GIzOXApK1pHISZBc2z
CAqL6kPWPbMqbVhwAY5ZP71LpYf7t/fK0NQgfpZz6BVsbwneSxOhKTIRoHl3jaQeQbrOAq3Sc0/f
cRRXNHYMgL8Wi1fKb2ue60mwpq0VuOiKmYm6lGavXDjcyioW3NsdJpmmhUkkc2N99I27fN5JITG7
EMR1lygROhCS2kI0ag0VfAFSoOijhBQep0qXYJ1rCip3THF5B6IysIpc/csW6+A+/IKKTNeuNRIS
+Wh+6Dfgv2TH15HFwwP/pS3KLU+gfefExjfmE3dna6Ja4bznNxJO9/9MB6wOdlmW5Z5oOBbiD/jt
3Rm6SXVLwS7XHhWv5YutPU6sj96nvQd9hgMCt+vJvgekEUORLOtLHNzIltw7vYYKMD2Vk0AUbAed
yT1SqarUGJAYnXsSHvLYpQty+Fnz6vtSfmI1T5I5+JEo3ywn6GsALF2cLpGe8hE7VAZF+Rmx4lgk
i713q9SF+mpkQw07GfbqpOg3YAxxgb1VBUgaMyHBLdAc5D9ZZx91C3p47TQZP6gfyc5kk9Y4n9Bu
8JVttr+A5m0sKhbE5EtKiZw2gyuCsfjj+xVkOc3pioJOI2mTT9UPWG4P3lUw38SmWlwXAHyy2eaN
XnVwjzc7EdWcoNSN7DVpzTPoobYO2sEEAtgb8paKvURQe/8kosdoFkN5osDtOTM6+QZgIEaN40pX
IMzWwu9aqtfvEIaLs1QMCHjOPNvFxrVt1+qvm4pIEv5oOaKIpMpUio9Qb68HHnnAsy6coftd/bM/
DNZ5R4wuPYQck8y+0mfRNG2ptIXZxbH4eOUFzNaz792HN0iZb12TBRRwzN31HEecm3epw6n27sIV
EIWxL1T/JqdoqAp+Ood+Clll/zHSAalmJVayJCtIQefFNJGsh65DYejnSOhpTlfiDV96t+Q+hfvY
HujOercVuhdpbPq53VRFXs1KNnl4QxbxvmEGneY8r9r1djx4/PloJdgfNNiKYGRmJsqlXVHGY+p0
WUW2qvd8Cf47L5W37OsMYXC8Me2Qerm4Bzr0ZOD0oRYc7Uq2/KwMV+hLUjXFnZq8Yl/4dDxtiBcJ
2NzSK1rgH2n1wmRSD8kB4fwaB74eG6M/thWUUhgamM54+lbziIs0148mMWgaTAO4dl4LFt0CWdTg
ZNc478V1Lj5RrUIvjytUa3ZKtymRIYO8ejO2osj5mxUruGHQipjSb02SdpwySR94jNMuSk9oHhtG
KXlbp006STTbP871oCA6/S/JInX58CbK253Fv6ovGmsDf4txwnTc/zbcWOomx+RlfGMs70coQYta
OClW7tDvn8I/ZmRX1RENqWvwgX+3JmIbhWl1FdPwgqSEgQZshGO2DnL3XroEnQC0EDxJKAImCQjh
jz4YGIlZNJw9b30owf0A5T+DvKsEN9xnhtLBFh2zKwLYBdAWMOcyjzjd1BLaN2dOfkzPR3bXwkRG
LNBUhWxyXCzHZYPNrIoc+ArYfKKoZqbRsgdBH1E/Kbs154jG9CJM+mHDHjnzsZ/gN9Jyzo3VkpNo
uGMHXw6UbrmScMNXkRJAUTSzz+vYgtYo7VCCEiq60Q10QGjuHyCs8WP2Q7goJjJLzzduXisND6DO
VYb8O+MFi+62298pTLM6++RvZdIBBwMfXL9Vof/Hm04Iy8cBLCu+Aq0v5ruJ48E7dnfkQC5dnuMA
OnnL6D5D7aGMhpY+Ls6PRguoGlhmqoR18vAjXRAHZp50Rpm37UUUjeTmeBclrUdrXwS2N599swEB
rIjwOcPdoomp1gtsdoc/hIWcpPT3y//xNkDTo1jCSbXD2A8HO+Rop78/guNRXHC2zSMUb95GvCa2
ecxWIo85cw6mhypexKHNdDPBOTBTPUkf/M9CIzfOw+eow+77N6H8d0ouC3z55FcH1cj8fk0RfjF8
nMPimA9qzUKFnF86bHg6HL/fbupF6HnYkc3zkeROWUKEJ6Hh4A8+1nwcb+s8DEieE7FgOw7H0ZIa
wkmhpat9GL5mIia68Bmiev2b0C5uba+08W4HpAu4rlsxQFhsre23N/LSFyH0FWKVJiUHClGUPMBK
t5rc2zVVFOn1dxrQY2rSJqWDCURpOtcEqSX4BiOpbT1CYmvaLPgrUVJvq0rDn5qqszUn1MCxoSVW
bxn5rJIrUfRCHmVcdFpeDEBYxO+X385rZj2xgze3J2gTpcxNmVRcg1/HwQy/YcawK7gM/l5p4DJC
b0vEmkBvH/6DGwRW58KQcuLh2ZVNBiqnDVygRQbb0vzF1AsDpjJsJQShAk+eE+WkjozRku3TIygL
Mm7vZVymrJImMnHivedhXJkM5HaDbo/LKRrp1NsfuyPlq0ibVGMHSpiBqXSRp7/fRb76jw2CScm5
IiJ7+kqhy+htpnl27iu8yhUcbCh9HT/FB/h/8uZLvXg6GNeKsjqr1MOGZ8b8YT+5O4pzp6YNMBvX
l+BobwHEIIufKHWOgLPrhL5HmMbYdsYjQSL/mGv0mKLWRwgsGz5Q8+UQcSY0oZ30UxAP+LGaDCwT
piJ+eSs4y+au7NVpxCJFISCO/S7X3gpbVWU2MQbtsPZnixyEGu1hC2NANqDRyGcixOfW3l4pxuKK
j9HWBEV/A1T31swDU8LRFI+wBAIAT5JaQngeQmgy4c/V42Beuqsn4GqY2mO5dcDR4ReBm6U50LfL
Lid/b7qzyo57ulYkGhEuW6MhxFgNKA13MktNtnitvXA8zSW2Tij0BohLg1+OtPaEUV5EMBaC1paQ
HIgDDmM76kGtU0wI51IsKr24wCMRnVlYr4hhiutjfRbpBOiUW9daBWmCUC0iVhzvgZ2C5emTwlw+
C7nbdDjY4KY1ZD2ZF3YlxaE7/L+bc1nddRfBitRnBR5FdwgzcJ87kkTcbViwEugvus7a4UaioFnE
1ug5EgpM2pXPuOUjukBn9sEeGO1cRsnqxNQvfELEf2+0/2AXo62cl5PoUP0se/vl0Ez6rC9SheRY
Wf4ASvbcflDPHgmCRMoXqdOUyw8eJypKTeMQGmJqfgkh9k6z2PELe4TkedDpFv/ZRrd1Ck6nC7QD
VBXpk7nRhkCYWmRzmnvgcl8htD3XdgTJpy6udW7ewH2RRULmKxwDMbY3yB8wgDi3O3qnaLVXhj7q
XaDp19gdo9WZFfvZJraL4ghyRfn8hEDQR7PMi+KLyALOFRMF8YVoGcgHgtBsLK7FdvPXykp+S723
aQMSdvsfrQX4t9IxBNrGaPiEgGCoXqhIdWnM+fgZuFYFllTMlileIYrFTtHiZ5Q5+cm8aRUyBGpX
b2xv8NbHnw0ai/9z3gdo9bpeQz7xYtVBDCoro/ONhcwi0EYGNMdZ+864mDudxUSMsnFMDK01rKeP
nmtNKee1vhZHaHkDJ13RPUK6qyS7X4f9aAmFsaxxtqb1bh2D+x/xWqtC+4tKkF4U+0FpWCtE4hF1
S5lGIUp0TdJ354uxzj+f8J5F133TYCOBZpcg1o4LnrpRffsKd+Hb5AhQXXnyLYrT6TQ3SIetsktr
AWV3XOAv82KnJn3SF0+9wfqEgQAdGKG6+cLTsZtFYo/DG4gops1szTOJlVdDjHQoVE4GomWmIhWi
Av4mrKh3DtKeZ/ozIg99056d8UkcbibJh3c6dplqyBeZsiqT+8HZIY3+T9p4zdynSPkxBhjJb30G
T4TIeT/YxRY628QeZGBEt+6l/tXGlTb5Jo0Ck1seGBKSjv+CBAqt8edTJIU8mWPlSXsIm3Ox4NBV
w9579YXund2vhfpYYytLuD565mjnCqSQqloupUvHHW+cQ9Y0nV1m1SRG/H8piwl74C/WzoTjF+mP
nlgwkNTgEBfnuhopLsHL9FA6k5zsp2J2qZp7c2PdwE++pbEk2cxNDudYN51Oq1J6h0Q3w3XI3WUf
BfW1MJch/KAaYlJnMzv1TRBfgQj/ElWfRWHxYvM9TC/yZW9zrJxYLuTFK4GSyZco7XHIg+asCtbZ
IkW/5pu0G5znz2ayNwbTHFbg/thK8wSW1eF9NnkQUyFlyarNqAvWImhWyTRhGde9UYIl4jwXlAcQ
0+KSUIoYk38nR3JS53W9hf6/OCNmkEhR6cTyiHn7MY8qLu+yzElDfl/tpp8pobyvP7B56QlS3DNQ
7866NJAIPK90fOPZFIR/Xuot8Nw5zK7H3MxUelWZbzE8NMCw7sGJjxNz7wutbByGXlDl5yBmqi+j
VXyJ7/aO6gPEtsJn8TgU37/DFAp7ftrR194EUihkno9EmTZeyTVZnqGXpoPU0TtDWzuWCI9KvLi0
ykosdYtNVdjaI8Q0S/fOXtDcA2NSfIHIH/5yH/n30PXIswLHNjOloOA8gjqRNq4ldKlMsakKU1gd
T6oSqKQc6fVV6iLyPrn5IaKL7sPtNFCnpPf47tBPZj59ndXsxDlY430jaEw30zPdQ+6zYS8wqgJ9
kBs5TTYzDSCekBkJekQ0p5z5TIoGSxGHs04yGz8KI07sZ9W3XEzeluznRYWuH+tGvIJmGmQemX5r
qicgBKAO2HmDgk7327TpNdZINqSsxkklvfTos7LstUZvrbK7JR/WgQoOTysKTBg9EPTuIfamFNnw
EEsxHihKR9neSqBRRDplt9dkvemLJctGIMn9D9h3JcBv+BWL+7w+0dg/m+yow059g7bP/xYzAIhM
sQruHLFZWpkZNpsKo2vwHx+GQ0BTWp0vPf70sSDe/N738PBB8ZB6EAQ9AVXf46DPp9jofImuo8OR
KOLQeS+gELRqu0AT/Vv0ixoFPBA9+SEAqsy2MtIR09yhLFbSfuBhyow6NsY2kngQyQ3kC0RD6joJ
z+3ut8y+rgJgi+ToFnyKQbaacAfF7XlbiAzXQbQDfghfUCHQvIn90rgDWXx6varIwmaVSjkQ+sgs
uH7D0mq7YwyMDPjKzGHSjZBTrjOH0XAJEsSizQVlRpPEa9Q47fO9ke7NCPxsSLvvoITSaeEMQBBt
2uF9xm+HOZlS/YHjMFF8srsbWN6FeTpaMA852kJjDaW9NrZfA49j0JRR2XZ4lgR4EqatOfztRBmy
hpG9CWwsGRzm5F8Aqa/4YcULG6U/uKewlQ4VYya7RCCj0TxDL3lNr5hj9SfmH7NCD1c33J/VLeom
Id7JI6hqra1RiNJL+8NfKR2lJG2CjbQBVBxnlMOYOc6uRHnwV5kf7Tqwd260FX4hrm9QlcLk7BQY
UDCCn/gEHxYbR/6pHXjGlAp2JgZOaMnE566E/wXQI5KAwi+Dgx3jVCnFdsKrZYrdWev79v7AP0um
jXXWXxddu5Q/AQCdYGBpdb/k79vbMaDZGzVoU/N7wKO2u7vRweLNI0BwKffzsjjs3E3H8UEv/ykp
p94oAcijgYuVxTbI7WIXmd5WSqTREkzhvJePahdq2jGIgQlzMVbMHBGPYqrHtW59w30jF30va8lS
bYb0rJBi4dzbDYDr/AdkdQhHqFUB1A3aiiONBVsFvSFxnB1HAlMamzHP58y29rOTFmJu+iW7xOe6
cZXYbnmhir9xT+tmE8nlQf+GcbRlf83CsxSyK62XRnWbOJqz1LVi/VTze7x61zH3zKzXRDFgYFVr
r3WpnE4XtlXS6urTsRKRb/j2MeMciTik2UZEz6hXc1JEQsH7Fh6eF1wlBeuZqXKQ9crSK0NCa6P4
qEIE3FTzK5Oyy3eRbnyViAObJ8KIj9yvtBvScuk8eA+kZWGrwRUZFibZb9Rz67MLlr9TyTm/8m0e
cKzVNWcZnPPnF1lYpunqSwsZm7IujA/bdEeibh/JKQUQcayTk/KKFgOEsbyG3KsiFE4dD1Uf926z
Me4dPhG980MTDRg8kzilKQFFDEZTFcQCax7nyhAfMjrOsP6GHEvnlOF8xtk6fHERk47oCKdP18L6
xMmWT27k3MEgGCbbJAYDodaTnuwfpz3c2Yz46b7dlxFrwUt3fJePEEQdsONxMC4aOXBdof4J5eGt
v6FN3V3/ud4E+MIpQqLo+vSuvgCU1zVCNM6IutGv3/c68LBRx1Pz/DAmzKvQr7zYTe5K11qA1nTP
t7SdMGbw0BThSTiOP0hO5MQyap/rhQ/PnbJ+T1pSywa4WKt4cTzGVULgMKLTemrBFiVUcX2Ala6F
NOslhWyY9gSmXe3cXtdRBwgUEWsUcTznGNMKi9qfNn5A9Eg9jkSyxkvfnH4ASs7lTbEyHqEaKMos
NKBwLVt7WTj9cObpIS5PEh8Vo3oXuNRtesJ+p0GEzEjmebP819QsCOaZhAppzDxzDMaHot4REc/O
VlO+GFKONrEuXYGTl9mmZOoDfdOyfOuyu43PmOHFhQ3C01asKlbfLE4eAWajuCsNpjX1xt+nKt2D
OMhuC+4jgbctQBcbT/ADf2Ur+Ek8cTqxvDWsCFrK4iuXxXKtK9lTjvv/g+V9kjYrI2qCCHKdfl4e
SYlzzUGVmx5CKUTnTTUVscGsy1gNwo1ArG1WRtA96kE+Ait7lN/iC9luar0oPcLZW/DiuCmmI2TT
Ig7Z1tVwqrTf/WCPAa7oRuHAGm+NjFK2s/NgNW4mMB7mBB9ChGZZGR5bAMksBPrN4JxwU8eqBU6A
SXfjjyFRTatbvvq8guzQ1X97iOwG2vQMCXPPZpQbjMABgh7H0ZFo98HFwQURFA64XeJW/9qtBQmR
ZQHd6cGhzrPdVtz34WrnBUxKQ7qTMISFoVjpg/9dLDbexGsEQZkVv695d/jGoCbF/7/aJV2TVPeW
OHAm23aAN2I6Z0dKy69TCEjc/wPt4FuMc6DJNeicdUleIfotD392r02sg1Xhpumb+z+5ik6gGlR1
QJ94u1+Czaj559UlcEf120CLnj9gwZJ4sVIxT+ecwfmpObq6HcWsI4vDhc3HKCw1VFW35tEAP1X7
VknwLJ/jq6IBKbj2ZzqvdJwGsIKswfSjw1zDjSXkRhN4xnAZW8v/D7JecA4iL05hgF22sdF5+LVX
eVl1L3h4aStPDIUvVWIMuCxNwwWkZINcZYHYi2Yb2lt3UObkNL2/Hm8hZWreh1yV8+8zVnPKWab5
H78LDQR7SGpgBNUgM2yZcjFqvDJ5Zj+dUz8uvOpcSO2hIz6BpxrkX04Rn5dcre3BkLsIID9YQgQK
XyNPy8PuqtwsZrGFGGQIk64lWrJ5bf4sWNdQftm/TDGcLfxh2KwytIPr6dcgMuDDxfYU9IO4ogzd
uDZReCfKU5z/ZAEnPP8rhULQUycnA3MBSlDYbu2xWhFWlb0tI2bNBRby6hqGzDcwHsMlQFCZCIah
O3l+TZg1fyFlwU3Z2U9e9zq7aDeOzRG5/D7iMU+VLJGuvTsGfa8n645We7GauA9KeFg1JHTGU4Ep
7nLXwMZDWAyJVVvqyY4cBNGK2I/EkGEC5BdayacW6zIk0gyEWhL9Z96NFXcpkYXPSA1WZy+u3HhW
/hUiERFRUNppajSyh+Dnt92HKN2c0SGYmUklbgdixVOH5KzXvKVGAdCkuDQiNDfarsgD6s00uVxE
n2lYAqAgC5enRIddbTt3cfh1eVQCltW3m7psO7FbcbYEyeLwNHbz2xZdfPgqIh6AwujBsVcKfk1K
mxbCJc3Q6nEB4ln0GeTfgbLIgzbP7SfQSkEwVcXCVGfl5YJFpsFSSCRaN64ZJ85B6vEhDOEQBp56
+gr1zyRwiGkTzDWUy6QRBSt8QfmGIW1t+LuDPWNBjziVDDKsX1Xq/7MUZzeyW4fjaXTsSVEgTSn4
rC2S1SC7SO4E9Z9AbJsqP4BTVHKG8SNEUO9O0J8Izqh9CFFcb55cyFNxd6ZYsHNTgA8sTOvupFCF
Hq2hv7KaZFgzon17GoYtXMRGkzk2NbqcSax6+5WYUStxvLNAsdjSl4XLL46BNHJWdP+2M7BXVWzr
AZDP0+k9wOlXlCj+UPiJnwawd/2DYiWWccDFHTvDBlqojPpg0ZKbM7FpaGpfWtShHK4S1WrqlPQL
6c4V8NI/XjxrlM/MPYIgu80gtT7AB6p1VCrSImVFGMTWo80xd15sZNWfzTyfHE9q2f+hq7GQRcQK
0VqzpRsGW3mkmlBTWozZ+pKOXgD9tcJPLsSk3RzGSJqNOFPC+fvs3+/4ShYSZddAbt53e5y/k4pZ
e9iq8ZHtO7OXHb4G2J/yd9ASxmrfKtGt4+UnGEOyUBevmTgK0hOJ5+CopkYHLua2mUlqiy8h7Bip
UcJsMy8HfwBLboNyIUL6rmESNNVqtou5pWyDkvxK7PZRkWrFjxowb1RSfUyRdz3cM1diYP7nhlLl
/tfmVaca3ffUcCNzzIZ0hWiiAtDU/Cj9rZJPegKFpRAPxboTRTo9TQrSL6FNHvfX7uN10r2Yo3oC
aUd1gIq6V8JOEAhxPp4ZoGNCCYFE6PrMH9sI6TI6nqlgKaEMekPc6ShAD9curHQQK1oetwcyahAz
W5GiGCdsAs5YXKdbsnsapqVFLcmqFwKKjGL5ERCHBQr6aV8gxqTB5pleX+tMmhLmmZvGNw95Dm0u
bq1gIvQGf382ToWGX1bcA5rt4Z98HWPnXIf5E9sfr4p/qM5e6EhUGvpzEEL0gv8F1dRk9zdEuLmw
lFv6Xwq8NsnM6r8QKwKN2IkJUlgFozpWaY8usRSn9C96QVguvC94iyqA/3maSfbqbxGRwv2+TIBZ
qQDEr9UpOjjmQxoYFIq35SF18zcPyqycHzF1LeDMbvWfxiwI7bXb36G4H93+RR0N7hdEYJHdSXH9
5s7axligeyfKdI0Yi0023wSwMqOKuRYdf0uctuEjyhKLuWcJ2OI6ZYLQ2JancwmGctm/i3dDVaAk
yR7LbGbQLw8QQREv1kQd8QIgLXGYGtWYKBbXNHgS9aHAEdZLQLqxtOnmjv2/SloMMvoQQUb0pyv5
2VffbrbyHfd5QozxtY7qXOFm1tSnySwBizIIh+cPj44Kj7RAbc8uilAbfaz1GzRuaTLTewWeIDXQ
Nj3Fq14nL4mo6i2wCTfJnKc9vA6BSsT3plAKmJHZ/vfISbsVw34wESG4/VCPJLDRI2XR5x1tDW1x
s5VlDUxETmNLYB6MkWaOrMFZtXZDeNh3iE7bz89l974p83OnX5q1BpJUIafhFmrZtzGWZmcFFPiF
LHdWkmlhU5Bq40VClHK1bmhkIVSc4B4ZA2xbIIjX4Mm/rzG0gMcJOUtUPOAHU3LLv2CGrTqZN08b
hBm01MExqbGUDHwrZfNRK2mLod+SM8srTFTISSFR9f/imXYneJEAny7FqegsWiHD/Czkc0XMxYxJ
n7CagXZf62LqjEM36QagPsroXMoUSwdTkS1zqJ3FgDCBhI5yYghLDM6A9zyezWQOeZS8zPjD6PeW
JRhLrYM7wo5nXiX458CnNo7X6xDMbufc/6AVjOMV588WkGDLvbTx/n/a7wPwN8iegq89109367Mw
x9R6eKiAadOKKj6obAv1YVJJs/uNmTRugS/mYhzC3Btr6mTplLT4p1MudROpJtnXKBrwiTArSW+o
e+G6r9W+4XXQBCIofIsZ3FMrxPhEZE0+orqFtn6QD1UfHyEW6sgDMmtIgZzeJOVJOfKvZ5DW0TOe
VT4q2QJCcV4s2fmr6tOXou/O+Bejl4y62l4WcbWN6C/CQKWPgnw5uom53YkKdFNEHuL5Mhgb6VZn
0p6chTx3WBTwcMnHb1IOEcRZ4qCXGsio9ntOF5Dk/cOTJbBBXuhOuqLVoBW10sDj2IBo1zCVnMCi
IKz7EGMaRmy5Yk0yYQnMDEC/wShfvTpHafDrtp0auhHNkzUkUPzWCRqRzg/wJXTjpknxWrJPLdgT
ksCrg2XUOIXVlRMyBlQi0JX6rlfgt1wRNeqhY2hu/lmoyhoC5AyCs0wQQCOsik/82g7t+VBrPGuO
qbfeyZQLbKwLgIiEWj8mrcfGMcLX2opD1R6zhtStQ8nzhppr9xZTP5ipWCrPznXS/HxLKLphVvak
VtKfL5p9eXhJdwMfuIVZ0YOePQPSj70u6tsSZ1AYn6kXRU37XoVltUWUW+kXPMAzMjn1NhQtvQ6g
wYMZuGxHErqhJ/9nO9HdtjTaSYMc+fZDG/XMiuWxq8C25clkvosf0l8JNoFRvcserQ75ouW2bAW0
qmIksmbAih6F/qEsBel0c57Oxrf+E+iGV0CvriyhcJUVPXHFBmXhHTNeUzpPv1m/cJdeM/4/9gBn
vJzzMba/cw5P6AmfdcGpQ1FGTeQE6RUjhGLRrijKTXJPYgOHq7Gofzqje94C9yMgcPOzrgosZA/m
Hid5U7C+0I70mlVP1VyBUTdZftqW0DFg5bKg+rF0qsnrhycYCascOi7R24ywWoYVAOBpHHz5aC1I
//Yg3AF5CrXpfcg6TECxudMs3vSF2cVuqfFDNmXKCYLPrm/jrcQu31f7lSZPevOCLX0L1zaC5c69
WLlBshD+S37z6x3nSPClamjRMgUcuePCShvMuuFmtRqESxYmf+Gy8POHWnoQSptXJ6KLfSfeAIP5
8tw1R9Z4fhHunYrepIXqncgpHzPMWFZ+HGiEsSJGnKf2K/J6BN6cM5iM6qce+vpHs9jZAiKYX5ts
ZETawjoaBrpDuBqV+14czM8D89lR2CS5khNXjkgSjNnagcabIY50z95oPZqjFFoCk1gBD22vKQwH
TVTzchbO/PyI3LefcIYPYYUc6i1XcMp24SVDtZKAiGLCKg2bqMErkrlkX3SfZ7gbXKsNdcBDSabu
rbiKMiX9V1FYwqrkPp51pRClMcqbx4+PDtX5WIhQ0Ku8y5/Qn2qCthJklUddMrdY4og30cfKYxn3
Gg3QYhNSnNBjw7dfYmOMQt6cBW1sZrHAoSu3W4ppwNB7Qx2F3htvqMLuEx8dvx/YFxbFJ2PxR0kC
d+WnoacDuwQt1FDQtxeyNoI6sLGRLIxRu7kiPtMeLeZzt077b6wG/2/FjBjgNLYgzxsOmz/xwPen
fGR+FXk39Kg2khwrU1ykCiN1knyVx6wVZOis9Hk+yxoHfKK0bS7ccLv7DiETP/Z6m5DLP2m78/jG
ehhGv/JreWHC2ZdYfBCZqB+y7/0Rlaa8hhY8F1Re1C1W3/iP7kd3RK95a7ny6UCtT5n4xGeUvq93
eTcyrEgTfvUQEYUIIZul93SNDr1A5kLhRGwFZlbvRDob4/L+j3TXeeLBrSHWXeFKemotkfG6HXWo
bF1dKnc51bg2vARm8RGNdUqCK+/P2FbvyKYoTJdJOOFlmukV2Y8B51dL9NaGLmYLGHUPzdI9/K0m
X62jF3GzDtd9RltI46unkOjwmfi0bUGMgHxRL9tucTYS/HyjkaAr2SWDDJ1XIuXiiaU8f4CikH+A
66rvyl34nYBhBOO174sQfj1V5C2uLlWZ3zEI2krY5SIN0Y/SZbuXp//g2lip/FWy3UANrwxx9zAr
LEDT6dyb7IPNxr9XDuQ2F2Z1jaF016aXf2bZrTQvhnD1iDJHyCnq/mCbNAGKlOjhgkdMWCRS+ZdQ
JZ034Z0AAO4YYymPONrkRUUy2NzjvJ0ZpxvGu0m03W7W0hFxzaqNu6lE8U/E8h36lPE743ZeuAZU
MEYr/2PTVojK6pCiK50LAlJUdn0VG0we1RQ6Dt3+Og41xM9axQgtlcIqNE7m/U8XYFLEIJ2Qc+Ll
1IRLan+H7owYz69ewZ55I86WkZb1uVgq3GVvWfQAj2SUrwFZ22KOBlyryO4et3xkcCX14Hbt14Rs
vs8KLV9qaxDXeUTwd5SbJKd9nHe+tTYHWX5qqZKqHXhOw5HRLf54ppKx/PBVnyBUmNbzJhWvzMG+
fmbKLIaNBwf2yR02gbdc7X09BnefXRiWGX5g7V6vGUcNSK50cvAcd5tUmh4O3+s3pYTIn9UqNcyJ
3mU8V0IwRkVjsqdBJCySnX2DjM5t9UFFSrGjA2/GncbIIkp5aTp/byGuo+XnU3ZrvxBOXw94BfJZ
72NMs7bSE8FujK0fBvoNpu3n0+6tV07TKS7MeDaEFDymJr3Fmm7ImBqRFgIxa4Wjuiby3mRr4tJK
5SzDQgX5ubmPt4WaPUaDaTR86SbD42l4F3Zc0ZbK7VKO9YRJ0myZKNBAPN4LmvY395bZKtDyGZKO
Lc/wjtM0dvuWVjVJNrd2Ki/UsfNRyLY3LeknOqEoPPhFEzEZx1ghcFcBKYLAVVjcthyUnflnXXVC
f20Ono3QCEtXmjPi+gm1PiFsLCjPhJXHhJutwaCpLDTLOK6dQ39BALYR+/NqAgV67NmL50w82U9F
xusWk65l8szGVHbqNGVht8ZX/DYUj+GDfecUQ4e8EF0dOSIcESAFmJZ+LZsmQx2VsdBH+N9JWx6r
A6AU4jf1Ha0Z4OUsBbDgvaWcfgw53ib7OvkHE5qXlc7tasdqOHVI5YSg/lrAr3LoZ4/MEFn8EGZg
4IzsPnqANiP77ydvDVKsU4YXLQ0We3FOr3d0x+C1WdBJL9PsbOYayfwsmybsxnww928+BjH1Yak6
T63z+jdM8QNjKDQYorQZMZLkj4sZMuWrTBQfTW15h6HrevV5Os0ACJfefQpGOkSt9RyytTIL2goE
rY4KjqdS+YOQbiQIC67wwdKWsymzA+NpOsdZ+rrOnfOO2sMnmN60nDqqvOh3VKxg+WoYj3P0WCvH
NbXqksNxElOoQRg8Zbt2xAtw0vv/0rqzk8iRU1gWNsh02flm0NW9FyPWrE1sEgEB7zzR+9JPXxMb
cG73zgsyQePz0WP8HyH4sOnqLGrFtSuSrrbL8nBHkpPeRosfbVp/lpukpX3hLHbSqaPbdm8rpuWU
OQ5Rt4gUbLqDIv2plkkbgkWSsY7/4IpUIm7zQNa7J2oykNPNsF/mVYWqezQPTou4I1kFTQhC6/L6
1pRFcTiAbHO2uWFqIQ16OM3TWkKcNmakQ26fB6Ch7Fg959DnEsKViYgvXHRPBKVQjsVLDNUB+DdA
vcTRfpaLRUZ9KBkbLVQfnA2GTUuatu3GYNOy2VGarNGofANCKNBpSOW73GvSmUCQF9T/8HMjYBCu
eBtZD/P3bXPWDQz8O8feO0hS383e1fUfRFj5uckxnYgl1VwQJL4uMGFgeUGpFJgidbo4EPVkfE1R
RbZWii9Ao50A9SOw+cgPVSEsaxwXu0X+Z8Wrj/brJyfqGMTEz9tu6c+jBov0qvz4fCahGeJuZFfu
mdscNeZPKrYTiWlgTn4edD0fZ0lOp82nkdiIqTyjxbZ0LO5odmzB4T9QYHDyZI7k4iWbVMFVWnyw
MX5L8fnVVQfybzNVL3vjfzwiah0jpUUm3xvjEYX/nHe04clqvU8phofXgWOG08HM7wXyltqoSZ7r
rT0tQJhrrCfWLh6GAvSm6gjhF8qOWxmRivHVCxNSfKGY0pKu97jNTNqxo+4gLtUvSAxxqQOs0n6a
vgOxOFa4I9FrEPcfZTuVvP9oiA6WjBxV1WT94kk3RH+7eMtYGvGuzy7En7os0B6K6pN0zreCmCPK
H3k8UTS1A5sRDBQ8WN5fCO1NTYvswyjRH8J84ChmujvFyw3TmpK2EDQzKWBW6OxvqhdKi/MzLQA7
NARyhAMpaLP7fAybF7bAIa5IStrsbNl0TsIP/x9E8Zballd1SLlmgfYW2Dvo067xXfzwPOc8jnpw
aHx2zufZBxE/UUXGrNkrIWda+tV/lU+LX9rJBtFm9Ub/BqPEcYXtAod4JRuRmNsvSritY/GBUpdb
yJA1bfBqlg3gvV1ZnxPyVms4t35qaqUfjJe/xqdibAWlDNM7F0dAijOOqLfvj2846Bmy9TdFr1WV
cx9wW/WUo27t1HOzbt+VORqCtQQvxwCYPS/2uZu45NnfBimjEk4lzjRsG3XY/yPGNu9skYxB/ZS5
1CO2Wzb1CKNpFJGI6A6vJeP//ThmOY0C3gNco0WVtAY7eH4elTEeNkynDhtzT80Dos+U69mkVZ6N
MziwkpC+ydPWGTUKnNt+ZrE0ZD8iGAeW8iYdlM7Nzgni1zEz8j9XB200McwjxIOj/yDfhGFjxZ+Y
1Px7skIuz0CnHaKz/KR+4sNzMYFwzeY4cwxBk8nPjrS6iHyzci4PHDiTU+54Slv8a4paMCO5NW+v
VumDM0ZXLTEJ4qJbockjPjoc8t4rKO1NFCSKbkXRNxIh4Gpb28Zjxyug4XWvRvRByE2H+PDDVoZi
IfihoDo67TjYMJthHry+o/0xqgSUILYnpI4E+kLpz9L20xeAMIpEzuvBK2Ns5MdRyCHOgW2XSPyN
g1GlVfVjsGU3uW/Na+ul3pjbplY9HTzqlJXEc6zbBnVyh/YD0kY9NKHu2nTSppWvEuasY5lmxOIP
HWqk4QtEsgbaKyu8rrtozzv1H2Atiba/YQAqlsz0BrUN6aJe2p7NpueeFZ3D9hRiWMSGqWnlyOAK
QG5aJblWAPFbo3KGFBwMilet2lcN0tgnhExtYx+oSBYPar0fKpTMp4O0zFE6qdhho7Q71MZ8l9+L
tebAt7hwLATZy3OP9lXgIR9/Y3JH9gEJpADnfmH1YMy3TIopnhJ5PlGE1tiwMpadi3C5ohOa7KQE
p9JHquiTX61VR63cAPdsAxjuzilDG5LfkqhHhOsn4oZQl1KfzNoPyNB1s+JEIcjF+TPYNtQnaiaQ
bRzRCDjOuyT2RrgS74fx/okkQ/hgDAQvSKbzt9ker/w50kgLghR2OLxXUH3NoXHtQ8j5CXVqzlh6
RJjD0WmVECLeqzSKee5p20ghxVVom7B0JKvTGs35eKPLipr+xx/QQoS0TEai3TVHl9SBY7vXpFfR
qnW8rKGeAxgOjy9KJiSZfdNDDdW08HCO7lrwpmfLzGzH88Q29FG4bwvqEm5VFko5IanYvA9DG5SD
wtN1SJB5EBkqe6or8MHD8csuTxY+6/W1Gvw14F5DQyDiLRwMNnB5jcuLTuALHIh9lNJoGgTvg/Mx
PNxQ3zQfTNVDWKe/Z2QjLt8gxHjLA2isB3D1QiAMwJiqZU3ARmq2a1bqJboWoR/0gj9yMF0t8DlD
+7fyvpgBR3iLY4hovOil8LYJ+H5Yf5Je6h0zZIxe23MCblhEl/RR8Tbz8dJqhNwaHMiejU11YHsb
ZIVB8/2ueJcDNRdM16j6EMtnY0AwtQNel9nX4W97Gmf3UreH50hoJzwzrFosJoWA87dStXyAq9Ek
9iUb3iGOz5j7j2Yyd2IeSQ66JxY8Y57V1WQV7/ROmu2M6SCSjyMzpEbezDhwCV3J2cj1N9rAbkQm
0QuYdt7z5eymCwgOjggDv/JGI0dJeyjhG9xpI40Rk3eoAENArk3dW1P6/gHOEViMpdq8wOeD1cKB
x2gEddB0DXmQ59Zk44H+JFswq+lh99igYfmvB41WLMLQ4muhontcbKTZPDggZzrKro1ipOg3Yc4D
q/Og3GgTK4zA8288K+RESR688vVRXayPnAbx08thKrbXE2Sr++wK4cEKqjdCJnO9EbnzWJXviBdd
EaP1+7yw6fOvjAZgHJhZqTRvTs+zqHkFh/g9W/4SEA+Gi1KqrN1VaR3qUqMBYV2OsRUuq5K7HLkL
QrG/V/dOKG0LdMAEyjjaQgAW2jA2pcHf7ornT58n6Zbb0wtikWNqpKsYOwu9mOY5lo6C/QOr7GXb
1aRdmaoNFJ2dtWPb21Uo4zO5zgaLRT1FJ6FoCbvmxL+BdyFT5X8mJXEre1GfMFytmKt8Oj62Mok/
gfYOsOaeb9SIPxyk0tKhaNz+rF2nzso+EruLcWcCugzlxfsnJz+cQdB5YhI7C1lvfmEUsqsS3OM1
o8gB0sJlY1ZN+m6KyV/2YTEc0uYdHyUmUPDH7YsRT/tY/bPK17Y1oJuQrQy8+Bm1urnPQ4yGIepT
Mwox7IUZaTtMhQnPFELwsZxWgLy1lub1ab0tG22wUFIcUasPBA3FAFk3oHbDm3b0cZKDs3DWhe0z
RA6DsPH06V/Xmq8RpXKWvSItpw8ml4jxec08hjBkcdvCouiaqPqfxHbWVevzOAcxx+k+k8qiSxFw
Q2c2l6p0GNo7sHof+G+Zkhc4TbfpflFD1LEdq26d73izWX3u1/kuktyE1ZPvYCLbfCu8of36RUL/
UVc/NsIpXZf/bVge/ZnT4DzA7vK17iWF/y6i7mJfeUq0Qx8OvVTYkHF85jx0FZrfswfBd31TcM8i
aSTN6xeEznldf6poI8Hfn3XzmmMGbIbVXYuwWbhg5eQR9a9iRtl/+vjuj50Nlk1DhInvjS2aTUUp
m9Y2i1AXSs+wZQ9i/TBM/EoyuyzwibUAd7ss38TxD6/zqx5F2PfqK4YyXYciJyb9MtxzrAN+wJAb
yW9b5bu/Fdz+DAIB+dfopPFG3ZfZEQsfUyXwPeW335G9j3a/Cgz0JelBMLFdoUYznA25dwQ0yc40
yVtkxgh2EjPIsFkeZw6rznozKDOgQVavHyzOJYwl+WOYN9w2IQ8hgbGQzveiAjqD7VCR8agMLhwV
M7OSOATQGGItv9I30hXyZ1zL/j8uVqFwUgPbzGHvZRj1uOU+UKoJ+c8VVHmBaDdQR3iQcCJpaZDm
YcEZyrDwLBlxR1XEqC8S5lI4hC5KqZqWL2ZUSyzW1+bP2TMcf6c/mM8hN3dUFX40guejNKlcjjTF
uOOsKGzbuhLSp4uXCp290JmiUvydigr93Ys5T21RO2OYbAvG5RHwHYRB7tEqy0+gojqFUNtL2/Qs
Ei1T1adoFJUF0GWfminvAPHXu6jnSl0CUa34/i+rNi1Ui4fvFVJ0h2RAvdKeWGq8VnL3X6jlvw4k
6E/dZ05KCLbLA71IFyH15UUV2tRMm8bHaJtAms01utHvxEgC8O/1eN3zMKZGGQGKaxUOZFh4nEzw
sV+52A19ML2qGQyAVQnJKIxQWa8D6P1kiuhao9Sqtlcmc7v6Dy7AzGyE2xbzl2PVhgTzMblT4F83
F8QU+39xOznm2Vo4fGe6VX8sDnYu83t/CCuaPsw3YHsI/bwk8yk45MthIzmztSRozgGsP+0Sjw29
CMNjIlBe13+rA+mk2aZVowmNOUnJHgL6N1hK/e/y6NmWqPEOk2gp9gt3G7wG6HKnKT3zsL2jZ5dr
yvFCz5Lt7m959os7SQ65cG+ChWcd3Vl7eJlDNeYvpOEAubDvDRr3fkFEGLXXEZ2uFPpUmWuQMXTq
7zUxEuRSiMZmMnZ5ZKP5m3sarYHYbgHGCkdhgxcvXWDUMcwlxiMRY7OwZ01Qy9HyfHozddf5mWM+
1pGJWTCR4yWyKWqwUYmi1DptUIdydXR+LyI0DmWd9x+BqJ01vRa9uud8QhDyczAA+I+7O+ZEeSct
xKxlcACtMggLSvJxNXiHII1KAyTRNgCOaATnLjxWly+vXy15OfSCFZeGKHn0szJD/UknRv/4HWav
Rq8kiy7HGgJ5E1nU4ipYCFSy81YpjIA36mWwsM+FElCgW+h0TODrOHcHyVY6qsJs5ijkdnWWgsjL
UQNQP5osXWrYLOGDqoqJeLKc/WKN8JUtdvqvnTNeAN/yF+vjIypkP/kShkXPWMoUc9kGWnds2Hwu
gOPrZ2fv9L+43rIBPcw066sMEy/OlZUsYXq0xqkLWiGSd5StgAqSBDB3Mzw1h8i4oqsjKKHrvMWR
stPRJY0noieK/qgQWKk7ufHTYayuywu1i7Z+T9UtKAUglcWwRdjv8DSkXHuhx6TSHjdvUVLHafaG
bPCxQKctdHM22Z43TgiQYQc1CdLKLLwsuNQbE5Sc608U/2/xrNoigpQqMuSay47ptliS+UjsF7+d
aiDBCFc7S1W+iFCfWAVQ1ux32KDB6Y5pAubdXjVyiEuWqOsP+Nq6uZ4v6KEwnBlbIUA9Iaci43d/
Oz3hrqwx+5xTlENdIhYMts/cu3ivjK2/OgJWDOsoi58/CbZZvsIquQ0W8s21O8XLp+DowQ7BNlDD
06Gb3veEUsdDZ7ohqHYdyplq6T7/1nW47gGEhg0ms1ggygz8xZ8ZtOTyeHrCr4B5jZT0cf0meDXY
wcbsmFdHRYVKV5T7Jeu1snkm6D+NRbM7qUQi5QgqWAPw4NDBEEzQPnN0aguIOxEeOI/wc8zcfEuP
gbJg1X6ySXmUPuOqUGv4DkZQmE2K+5IgIaYzlieEQ4Ceb0Z3EGNHw1DqyPBqwURiDLLOWK/tM870
CDQl3s/hsc1GdybSY1nPrLaIuZ4buKPTmYFJGTIQoGzKqnIVsMRA8BkHntTAc0uVyyou3U4imMg7
ArJi2zaPfRUNwpSx76L1SleE79nAA7f3Q2yIR5JVD9T8ax4KpEzakvOfBShs9BVVUC21WRRnFy7v
TBwPmgVPEFIXioi52wyo01aAGPyy2PGl2VuKGxernIyQOtDp0Vc5xH0Dz8Ckheu/eebrUOM7lGxM
+MW5e3p1qHfJvi0LQPrYpS/GesczvAM75GN+DREImhEgHxJ35XQFoob7aGeY70J2asjVRCwWPVTf
WnKGW86rNAeuWQog7tLZuaFgCbqRun8/apqBicyB3vlHLZ28/gHaAXF3O/NIAEXQUTMitnOF6LTa
6+Kk6F+yYTmwRiDBVffqR+2qA+oXN9/9TkVrvCTc/sy56pkeRAqp0ABJGi0o8hzpLc9iIPnhtSL3
VlyGcZ3ciECJg+u6lYGFEoUJPFord9DUKgZh4aasKOdRuxXD6cFxb5Q61jWccbewSFjmTdq8+eFh
ReUm83wO5209uODpLxuLgKp1fujkOks+9DN2RqSZu8qHmCJJyJcOrekqPqPctBgYSOeRsIHuBX34
AvL8JX8w2UaTJ4t7LFWhmbwAwmQtz1GZqxQ4Bs5Nxzr6FPB8hh5aZ32yU6tFD3CaMXiEd2d5gUtV
mMvPlvA3HLlB0cTpECSU0p3p15U+OwAUViswy3Yf64mGRfjjYgjuZN13RYusoo1zuRsDsng24f52
2JNDj/1hmQ5a/BkySO06kjCB9rOtNXVVS06jWpLBG8+PSoU1nKjwZbKgYpd5BV/4I8De29HUQV0W
S/HH9tw4+MvdpE3DJRohzZh60DOdlopQXOPdjxTyQSP9y+ChxABYILleujX3ae9cODsY2CGeBo1W
NeHrVdx2YJ3Eb5tSoL+dJhG0/OZ1ZiD3JTXp7Kzxme8rzx/yG5w26pID5zM43C59UzVbcq4aR5H5
X5P7HlLV2Uk4vpCiSB+aOPYunJrkLk0obsOLPiZhG05mwIEfSeDzkoJxyVroUv/x6sOsFvYoJXnp
GRiQzmrr7PleOtz7L10pQnGZnLQMwsJxNQP3kXRDM4Eb9V3+5t6t4CXq3bTeFug396WdEGt6dh8f
uUXdOifCOtVIRwxLVYA0wfxq4xIeQFxRye+kH8IiYmE98Xmz99vChOwnCs+1c09Zd3oUgIOVZHyw
/FeYDW0GxfiENWiPfT17h2xtfD7slv+ozZEslkpEwpeBgcQLjta7Hzqj9rh3bLGJ2HAkvrDzfsfJ
bMR42pbrKocSZ3i3pwaL9EVodOIThFTGcRLC+oZuHi57tbDqQpoHzGIOT69OUNQeiyudXr4pGqyv
jfX91Hfa9/C6cbnEik0Xgkob2fbeb2mB9iNnpd1certg/qNTfOXMrjP1U14IuNWJ6F2v5CwSkeT6
08aQZioIgOphUfJ6GfeULgxQLQonw4UjfF1zz57AXqac1dPCTNhUuAJMPniIjuztCg/oWmk5PXKA
XRNXdtry5GZVtZ35j5vds6uoCZiwUbIB0W1/mPrqA6i7Y3bOKLklk2BEj6mZ6+X2s86B2zCDELrv
q9Bo0fp0J6yUsAO+F2qQpII/oN7dqBEr2RDTXRFCRbKHOY0evZzdf4U0GgoAX8bGM1e7AbHbv5w7
Q9IvY/uQtJJfzewFxjtb+jkKY7b4CFlYIjbNDS7KLrXdJkQ4usud0MsU3FeRwePwhaijYkS2+beY
IU5RqpsVZLukjnbuFETQSAgFTimiT08eaI0uNGOjwSuEGQpFSFBC77iT4m8lcmFZYrrwPqSUsRx4
SRpquyvue6kyC86/gFaaWndICN5THJHgJAUNrykeKgEQx0fWN7I8I9L0v3Kssc1Gf9eafF5GKPBT
PV1Fs7T2hVJnFX4a1YaeZgkfFKKe1EQWVyhO6mJwXP0scwIqJDSsoxiGK2Qma1VHcJaQf6gcINVA
mxHXR0aZNUmXY/zKOQIIelXuPJ71ZZFr/3mhge015IOTU624wEc4hJxOA1Z7TU2+NQPgpYEa9y7B
CB/9Bcx66NhPS1zJ7zTZ+yMDVMNST7WIjUilaXnYKqzYJyzxKM/4B81PY6d3R3omGd2KXhzynQhf
JdGOZ/cpaSTxjRgf7n7ipIWDyIrmxWdTaAWOv12uWNkhtgEMUg/Rc/zDsxzPhOZbYfUCZ7UcI3oy
YMS4h3By6bvUDvGp5+oK9GAcY4UkpN5oSQqLx3DYdwvMRTHVi+CNvHseV2DBH7d9JNdgUZt5Vg2r
HBOOszwOZd3vpS/JSVpS3ZCWL0c2F1aFDyFfSfBU1zj/Em7DHCPV5hV5t9H1ChAjKnVEDCieesp6
4BGhzvWtgPD2u2d4wyLwJAe43gpj8XvBugGMYVBoJrSYik2i3vX11bzwBMOW0K8bBvK3x/XAeAEH
uVzaV3JDS5ki7dYGkClauXjb7s+cOJpkTWtEM34KjIaOdg8sYUp7wCxV3BMwcqGmM/Rt9YfLm/kI
eyxURAu8FBobM204li8lTEZGi8TcEwxHFSi1I4h8ki7/wJesi0/Vchqw3gROQXvYm4EzWAFY9Y3B
9tTfbLuSA2v47YA5HiqKElqzUVxKSsGJPNKGFDDzBK93+gioAP+R0Dj/JMLqD54INCkjfebCdiAe
663d9Mshtrq/uX42zT/ufSFuYfj6HYeGU665M1tZEKBgI1yk0qXhXdYPMgzF1O3vhwV3cq4aw7dI
Yy0IknEtkNPriMZn3uigo5M1re0xWMji+xoJMwtGb0OaDGNLDOW9boofpStnDo1NW/EQ3xOoZ989
rGa9CJz2NL0Dwk1xeSLqn+tQzJutNqVOfQBPch4g0UWpdNILR23wunJklhcZ1eSwzqJpFAQowSBw
p7XsyAr++YbKKR/1i6FHGS1jSzr4MIgCV8p6S9K6zqje+07/ypQf7muh50qltn2b8TlDxxVHmsbS
vmzEe151a7P3L6WqeW+CYRlZgISxJ+NxSPKEnKPXkOEoN9bE4ec7lp1sz7U8GCfiVQaDrWHfg0lc
5WzG0teEDQouDIsc8OudJWse4tSqMse1gnr9+z19Q+1li2Nlr2OCKAHBqVkLtRM7v20i0TSGMHfw
L1CUfoPXZ18Zypr/7aOeAryLkluyzrS98xlNOY2qniuxZk7mw71FwqKvrEzuaozvPno6vrQ5R5d/
fjVY4enallfPNn5asTGOyxJAx7yUx6i59qP9t5ZYgOnfFi6IMAls3CYFW638z9hHSBoymR3boZE5
LzRDerHqwTWtRLx3MLyBRwoFrDj8M6b799NYaKnf1wv6XhBZFt14LKbu6MTIxqilzK5WYLu8+v10
EYBJSRi1Kh9jVAqhkZX7ohNkl9HLv92lPFVP6W4QYEjxeOca0YwLdetlxRyWlEXpiV+UatrLQPkm
1/Hs5hJtSQcv2ZPdMup5I9dzmvbe5d/2pHZ4IJkS/pZICFjEpoUO3+/Qqqkbj2XATgzuUHw93Lgi
1RVWZ23veKAoYmpssN2LHXHH7UlCigysc0SPzmSgl0h8ea8kmIwrLYPr73iK4iU9EfbLuqiiMFjW
/i5h1HpJVcTUuwkjnn+XpBsB9VzqpghN6tPoPC0Pb+pMcnzUHc30lYYzILbuu+2XCrAx81jKWhxv
8xVRMJ2G5xSzGr4nXkrXxoceylqGe7FtK9a1HyYtw2x22CWlRVkVYVtzwFDTH7iBupmYHf+nyfYD
8YNg5CgJMrAh5pfjB0j1eSQE65Wab4hMz5ykBCfQ96OEBoYETJbkNInwDEQPptgzEYpClzTb7hnj
BaWJvhaa5MaBpITck1Wl/GUIFFi8e6n6sBBV33HeswlOdhu6FMQW+2uh6XCcAk/LzBCuwKip4G1w
1z4ROqO0ttYds53dc4N/wf72EI0AjEvCpEBEOadIdMh6WdWRya6iYG1m5K8iK3YjfnzfrRHzp3bI
K3QjIgJrT0dQJjaf3yCkA307KkUC4L3ZTwTLXrTY0u3FDo4Nd6/dZggSJZKqNCxUO4/Q8ACCGdic
9R3iodUGuSn1J6+NWRCALyp33JVNAJKPgKQdVebNtYtnQsKMm32QVdnNs1thrhOzwP0JIG1J34Mn
qEyIjCemw5FGx/+qnmArImcAsWxQVW4Ci1CcDL94NtibgE1QZXTiRz+jmePeGKcXvVDu1ctQVQ9x
JhFpYbSuldbYqOCeT+dih4xm/R67SUMvnsxjZzu1wYV4M1JYiPhuPrRfWR+6YHjRI6i6027V7Phl
j9eT4SpOoihPMSRa3zmnUZ2YmA9I8tr0+j2zSNVpE3FcwjTeqDx46ha13ULInPpPWocv2Q/pUYM7
OIxtT92lzC42pQAfoEXU2Gvyhl7JbEwrz2R2cYOYiRNLsMzMCNBsa4JGAnWzJ7dbDj84cRuhSOe7
3BAEWwyyVmNfP23bwEee/Rk3ny7Km3x6GZDSonCud0ZnAWJ2TBFByyqnUrbeIa5TM7udA3SiCPDY
dxToFE8AYBeXnpNkozYHfs0vXyHT0GZBEQ6crgPKF4yy3SToerg0IXRJ2X6i6+f5XXVQIhlYYS/W
PMlARe7lD1ka8fCqStX5X85gPS2i1jKg+lKq50w38w9x203Ax36wadiC8qw1745Y0mBROKMp8Seb
dQtITdjV9Q5dd/KS/vktJzbHpmRKewPw6ihPT8h9DzVzhlbmhUpA3GtqVjf92lOarPlb5g6vqSwS
TzWlaLSdEwqHt+Qt1Tpdo9S4nrRj1GZs6d2JlSK5wNfzQRseYIgzVAndJmicM3hizmC2rF3wS210
L6tnNxF3OTPs2hn+mLRrfUhZ4P7rRJHnKjbMpps7K2UvuuuqvZdZikxwzOt5ytR1mKTypvDicgNW
CzAhxg/4sRjSKFXPsKygbmTbk/17Dm9oRqVbD9f3+cDQGI4oc2zyNkcMdTg0femz130d2nOj6CVn
phG50K5nL0w/4llwW8heScO1OgAHmaxE5F90/zVGY2bfB1sMstobbAgaWxTI/bXQU1qe0p1aNmWg
ePnCVosa1kNxGNrV/vmd+rJhl1FcZu4ippaoEZPUdYj2ZxWBYqiHWo7IF99rv6XJ+oBnD5sBh5yG
ET7+A8mXlJCqQaC+HjqJzJ4WcgAJYXcJoLDv6vQFKxr59N/q4H7aFRIOosL6EFLqByFZmHn9YCGK
nGXxvPpZaqPHoMan6d0JpVVWtDpx5WJYr/juuth6jV+QPSJHQMD94vf8CSzKe24E8wMewf0XxeaS
q7yG+RdOyOFSuo/hRBQwYNbui1k0xFyjwZFGAZbB5QQJPboVUIrqbJ3zWQX6BhlkOdNQgovav08+
OVeujY0oVy+XxGSeT2FFYXw5QgspNlg0CqvWWzYWpZjiGoBsz9fjMvXaySQu2rjMwfn60LFKIQcW
m4NSchg20S9SA0XcbqzQu1vLm9o/jBOn3dj2TR0TN/C9FW99bkmA6GP0CAgnBzi/rpmIyRDSOCQb
h5nSqFO6JN8enVQlhCs5xA+vmNGrCCkFdXstNHvTJfAinQqhRhFJJfxrC2wFEFNZ00v6fcL+BOZX
X03/vi2Dergj69lEct0tKN5zBT81OF66sNOEmpn9PQx46Di87MN7icvcLJ6lbsWSEGMOdSHhlvOI
YQn3+12D0dsfAm64FUwldfwghlZUmABpycmwTaar2DEnok2ku0olVt7LarE7HPrOAy0U7gqOChZ7
vJw21Qv4V8hA0gNa8ZrkNLbSKhVaCo8TN7KKB+WyRoxtonfaqsP3gxW7Dl/Lox2o3q1hVf+cMgyI
yBRKy+LH1AeLhTOzKGo68E/FI/ONgfRLsQnyfqZkXp4f0Ldd6TNBqPehZR9z29fHpnRd2WBSShp8
JGv9hjil40ITxMtHbJgmNjWtGlqqQXXBjaZKKkKwbOp36o6gjuGMlBrwCMjpcQDFj1Zkh6FAmB4n
5Lfa6xziAeLl0elB6ElCzrvNsnA5yOd2W0T2D8190k+K2AYnyQvTATsI0/HWaCPjs/SM6S/apGW2
VU6kwWZBYjAoH8TZ1/TurGNFHuoQZDfsSgbZjHEcvZConhbfwAs4RZb2oXZZGFRo43QniUAZ9KU1
wafkfDbJsgq/cgEj+y4nxYaOcwx/xTlYU8ekRt4EgzmYCGQxmrSlcEXrIpmYYi1ZRw892py4mhKt
qMG6RSXHx8yS88qWXvKmathb1tSp/rGSN6OSEZpfVgDty2Rlvm3aoqg3PIl/g7nYW/ltF8H8POFn
EXzX/y/ODYxwBNPQ1ERVeemkkAzha3jJiahuoc81BUj8Br0DmgsZM1muYhKwne8AFS7pRlGCAKm3
ZFsZL8osZbRs6iKfLZvs8/GT8zyhIgOtelFchaDykEzLiXEFlYkR0QaZULhEuW5m4SsCTQCOEry9
oPf9x35aZ8EMwOm7QMppWbPCqim+HNuYSGjnPBQrFtcrLmBew+FN+6A7Z3Wdq0cjiXB9IXv0He+Y
ZxNbFKWqI3XB7v0RApR1RdCLwVjlJmPByrxmkIqnKc92VyYGlEBzrHmIFNsF8JZeacBe9QA87vhp
J/yIZpbZuaKr7LII40U/BxGrpQhR84GyRAS3i8+4vYSlItNZXR+PnDQJEukWCzBAkTyWQwff/Bv8
+OPefKjkNIcFAYJdL4IIYvzPyaTif4xKo8unAtSJ03ZjdxpYXFYd4fXWABLkN6eX7v/8MgLOeaxp
5ZG0b8Ih7EUxbUPmKf+iZwo0uiYhZiIMgdHS9H6VNeLq8+xu21eflzxB3CUc6yGOp2UxK5qQNBDf
YyvSpgaehSkOqXeR5E9ghTAsBEEagEDB9H8WNmmqC7L1iTmIMJVFSyvjLYKx/sikfzOrQuO8lenM
UStuK5PPqXsm5lEeBtm88E8RVdItr4OsWkcYyMnECh7Au/yN7AMKBQR+TEaOebDGpBnYUcTQRCaC
GKf3px10yABsi8I08poPlhmZv9NNguWw8a8l5xnde2k7NzNuHYa/wUO93gu+U9lz0Gk40dm2qOgF
8kPZBJj6HSO8MLGCOdkCQxeb3IMFdpZBatI4u3Hmt785nxYS0RBWcU+qRg2J6Y/pkwMGXXB+o48e
QVnzhiytMxeWtSHe6YKpuBhlCd/4mz8xA7xn2u35w1h3aBe2i4K3fStGoEBdQG/mNOhG615oTElZ
0Q/w+eQds9JgbAaVfqNxm3Fx+5G5/ygK/aDTvCJuxua/9ibA2wsPexgsEt3A3VFbB71E4mq6fCxr
sKi65YOPE9wK5CJf2I3Av6sffQdZT3IBYoZtZJewOAEVAYJuRGcZLZ4lAHAMEclD6Y8BUZUH1mN3
MM/RzwSVJaSu+n2mRg4FCsTkbO8tSEXevKiA8Q+pR5dNFsHSSSUz9a+BZLZE8aHFXMClN56p38iY
pOqD/eYTAwpNmRLzYWBd7WKHNpG+e/YhorfM6LwoW7v4sWX1tkrSRfQjm7afBpHCXXPI2/M2uYpl
88AuU98PMV1vEL24LCApaqI5BbaNRGyP5uakqbvHT7NpzDkY6vNj0tPJFHJ7Az8bhUdQ53jAOjeS
a56e9W8MYQR0FIsMbHuOevZR1jSwRazrIfaXYxrNNrz8NsotCI13Dz82s0d70ZTxDuE69WAX50fW
fmSRtU+rGb9m/qMt2rrNxXmv7ynjMHqXXIy0ypDqlyHpxXMI4N2+o4H7MAk2khF2juUYcNZLRGnb
R4Mbc99hsIIOREgdTM8tEAnBxrWeS22t0M3hiTOx3iLLzt/SUrewjdOBijKq2MC+MYjGNkbOzS3l
rhJ2TDjre9yDfO7Y3V71GbLoMtjPi5I76/ltpswfYzwA9uEAFs99A2Tlnj0bNlU2+CGsexPr6o6l
9t2Dm1TfBqP/vhafM/KT57nzSdTQmNqvuELPCz7O5xE64Kdgq4rDHuzhdD7/guX4xpgSrJHzRpMI
y/IZiJZivnONaTWOLdDaz4AUd654ZjxyVYScAnVjHFEtGa4ivIHUlcsRumCLM/czmCZvKAnqOGrJ
/QBDFELztKi4WbIrrkvDlPF7MHnjidxwOFhq4DWYv3eXrph/CTxNMUhC8cYcBaPMPmSq4VmKsqWu
R/w18xyMjT+d66pbTKo28K4TwGQBmKSzUicFK6xETkRg3oX0+S3xsyhugTkqxLNN+H3kzAdogYyM
PUxGqp4apV0A34S3GTsWlm72GWxjBopxnz/kuBRPbT9k5MXalDxaxocKq6BZC2mMkMBrFfeSj83L
Iw0vp9rZgNmI/2ApgnO6ijCDWP96LK7AocWuCakz50V7oNpWYkHnk6BLeiizvnwD/2f6S6ABBiCb
DeBPmwVaxz2LwEAXFADKboHgChD8ppDe77B505wDGV5KN5ZTJSMaCpv+4RsMHyz5kHOAneBhJ7NA
S7BILlORN7QrD19K8qcvlzFGiRqYSMhi4ee3U5XrudZOEB0hOywidLkrZONcgPmkTRIRuyCeUC7h
bhWq9Sm5MfTCx96cfq5QX66S51YGgXJmjaD+KUqfHCb8v/JEwHE+4lit0MmueF+DiTMv2RKml8Si
z10F1AsaWTvssQVR0RIXith1zGjcGlymoRsctqoAF+LgTzl8zlWOk5c4BoN343r0/m3/nLN0jpaz
6qFuyFMQP5qWOcBVk/f3qfRZ+ZHWASHABT9WVTouS7xpb/kjq6yU6GHK2gU30cGpc67FR3kQhS35
vesVRKBzeG/pAiuqhoTOIJI5YrJvcWtszSjTrx5EF+S0jnSJJERNfzOU4Ay1WxqUV08vbYL7xgvz
4QuMXCogfOO2wnfK9GslJtBpief/SDT77hyWvE/rHXmmCSA5kjbTuav7gUjCh/jsZ5m7HPuFAwCr
NgmXlh4yI1MiL0Epx6nHzQMB2CZdt/NQEY5lVeC8W4WOR7qr4FHaJ9f+tdtAKPwK9FPUC4pK4GC1
+Lj1juO5w0xSPoLAUNmNbbckNHS+nBgBp0QRXxAY5WdPujmdqiLEZl0b0KlimItkDtTuxvimWU6E
DsROWIRJH5AjcpCI2EB0XHWfGdUONBQdPFsub4mrkDIQ21nIBN+cS6NdfMPm8goEYlh1N8jEFPKy
rsMNzJFXJLNo52lDJI2wP0WLeytJ79HFxxeFx1OZ1jW5ZLF080gNZRHsfNwa5a0uPB8+JO0chPbX
joPxoeFdyreo5Un5Bseuyr67qwzitB4gyItVaaE2HUCJ/aIngYAWAj6m6Rn0tcBVp/5V8LWgwh/4
GvDGyaFIeeOWPfOELObTPsYr7Eq3KsXqudZVAF4J99iAduj3u0+g0Risd6tst6btDJpz32f/h1BD
QhJa9H46AY+hHGHfh+eMAHIf6crxk8aQKw5ZT5WcgIKrSKWhJ1vy4ZMplS4/i833WsswRFiqPM9/
q38qC91wl8yiSVawRNSC2YCeiLzynFd7HPXZImZlGA+IcorrJjrT6kFUIPs1yXke135uO0tPAa3X
A5pSzX6TElTrWisAdk3JHSQMOrS4Ye1Teu67j7f3g139STx7lkyiLc6WzbwR6UJsXk32LGehJzaX
NoqM6Fihe/u/mqhhZY0L1vC1rljjAuiefY5aOpgLAXbwaJQUcgX3BoTnXnCnVw3XgtCOVI0lUXqN
cbs8do2vRdbHzjOG8DWSZ+la+3pUfDHauzmGUy2x91VL4VxJQuPis1s/NiqX2unJYuwdBCOQnwxR
J3c9Hl9FlKY8+90sDR4WZyT6XMaEivHyilFTuauH+6u0K/3YHAA7S8quVb6NfPxejfDRobRwcHPO
rYg966UBMgiD+aBKk7M9eLg0bFp+ONWDJkJzInWJG6Fa4XsNCKKUKyCinkFDGsZgwjrqPCqQFlgF
Wxqg5puqRUs1kWeyhfm4+bNozZUKGfPs3wGfbdYFd+Jq0gZ+kMiqAm+QBqi9MdVqAJlbYAxlGSi6
4fP/17VjdZoi9zJfiUCKO9733lGO0zMHDS0TadTyW6PegJPGtzYjX158+SJkysSE92ogqAEq2COV
KNt2S1vtEjg8zU7qEFlpIhT395daOlURosqSEd6gA1/WGWDX+7tauUzldIAMJToJHHplltyBo6Ia
blFh7Ml15zdxJth7nYZmB5TT4/s9UBTKHrVGALJBdp/Lxb8fAEurDRf84G1dFSNBg3oE3a1BilaD
xOuiHnnLlEG1g5U0pGuVXFo1hYA/WRhJf5euAh1zBOzP/cN2tzwKOFYuQLVpMw1V9Ax9ZA3RPANp
T6/bY+onZBdZI/wsbtm0Dk2D3GsIg8rg+OdOlNSGh0cueLAtWtUYc84ViXU4a0+aTbEP1czRaezP
KsR/y6bDV6NHZzfWfJvSZ08c9XY043ks9weUb85iByBbOTbYtnDNBekd4Fb7rILudNs1BMzX0MRL
D5j+KJqk78vadoQfFG32UmHQzZqd+bzNI5DDNtjmzgFAw9P7WjpZOXiUZSRIPD7fYNk19YFnNhx+
DwROK2MFLdsTVPt7xTuDn2sFUP5+PAbGL+AY8vGSd+/iOk7NAFe+tR5wVSbWxtxpcgSbP9OjYErY
wCnBiczO7Bh/IgH+zvDORBLAfyUC6dc3Y+MpNOrb7qCrmRysdRroKLwaMK5G72a0wc0VOh+toyZ4
KJTzCLRvGKq7ulcZ4YI1pGKcUCuiw3mIJvVpRHTDibAkAr+urqZo0GgA+jJAqFXFSS/wg8YYfYJb
ADu2ecQBZF7ZwYusfWeSx4k0sTEgHL/7lj3J9VXeXEF1BFsOcmn6iO4XC5JnmKvYoHLw0DwlOe6M
pNbrKYXnlHLP3uZ+a3Zl3x2d6G8g6eVwwp/ZHVryLRiEeDJmdftw0ccdT4atysuHzCUCz61BBFVH
ZNlGb+wTlZFTTBmTuopKHa68H5h+6x8aDicLolslkOFhCDu0WJI0Cq04O+ymU+z+7a9o3DvTnX+M
iQVjwxP7a5rI6Y5ldWjV6f3mpGXV4UwcEH7hzdmdK4Aj7AibQCYgd9/+JAyzRihQDxUbo2Ymx3Sn
011bzMFqsob9X/c7/5lS859YjhvUH24cNRHmFNGiqcXeoNtiYjjUItQEWO58eyYkQV+qtllVFnBl
dznhI+7jgxqnonipSmApvoc2XxWdZqpT+aDRWY1uMFuPLaD7c7DlVGOEDRVp+alnXj6g0sevIBYB
oigjV/+yuEwoNp4XEGLhlv0AC0vUpztqVKKw3h2m/7G4vpX6D6dQdVwp92/1nOIfZUv28MVv8Y4P
eI5UnneTy0cyd4OCrUidfj5xEBT050bJylIrj0bt+MXCreVHDlydW2M+PBdNC/qzS4LJYFDP5jvK
Eq8DugdKZjsXMyF3+1UxqTpnyeG/iGl9N8+m1eL3WXrT6iFnUNrJUun6n49Yz2eOD6NmU6STkRZj
Hl8AJE+4IWcVyT/EvOG+7AmlZ8pC5Th8B8Gr+3VaN9chbPsKLromfGRmOaF1sKdTX/qNmZbelZRa
1/KxWhtwY48ocl7BbXgkWssa6IRKVpjfz1XHK2HId8e5xuUuLmh4mJfnXVl8GacNhEK/fRkg6OFW
U93RtfzLX3OnAaCaz1/sav3k6usrBY4/IExi7To4e9hRZTghfPUpRkwJKDAO8eRZX/Qk3MF2agW4
SNAHdPxenKCeDNfoD/JGnQjN14HQJsT56lawQ6tygy3/b+o46cvTLEhOFpUvgvB8aQ1phyup1GIT
OWuctnXODFVeCm12Pev6gHPuDamD6K/dpRIQ889ypfiNZziBCEjTEzJ9gwDFfvKIuuq176KDI3xV
ZszCLEitfQiBZhgAABiLMsgQQb3ug0ayK1Kt2eKUilUnpKh4U4MpVtvtdtuyl6Sr5MKk3na84Zri
PxJ0NQzR1dPbGBRqhJpYMpvebfUULOH+mlPFUGSE9t13a78PADOrZHmZ65FV3/J7wmB+wakMh1+H
xLSX9/RbuzkDbS0CTqkFYOt8QnzvkGqMEbV9DhRsqvoH+g10Bu3PAuF9Xr0K5MMoOkdOnCqp2Wvw
9i3tMiLSqi6cAk+XSEndKZpAQKvVtBG5dSePmI6KP96Yr2uhd28iI2oUzp7BEP5nxMvDwlPzeSlo
7+XjjYBs+RxgFuIHSgo34rLc+v9dLKdzLUUldA9X/iaVfDekJjUfzezku2US+upHQHW8+NWyCouv
uAYQydUGQoBdSs+CPjQbRHcwAaFmYaVMe1+31IAq6qSOZNX9TH93bga4IIPLr9e525i7UHsO2UbQ
K/ba7pTbSHy95qVX672FdPUXhYOnX3n55g36rOMKzO9GwdYxtl82pfoGA9UnoalRV4CH6XTvXunZ
cWONxE+C6j5Ezxdfq94AJw1tTlFyim1AhhZX69Vmbo4JoB2UsEhdqt2TfDyl0OlrcMadq8HSl1dk
Dq/w7gLlJnZsbkncStyHMvFNjfr8Zb0/5Jtkq33DNymsl78XON2iIF0G/fgTELl+iNSejb6eKXRa
YsSzJPIXRRjYkvF11LtRXjYgjJi7jWj3ockvhg/8o1oXnNrZV4C40lFBJpKp8QivRpd/Mrd6DUO8
z0p861QyNnElnJumIZPFuNkBushyp6DncqoftfGBuYF+jQLWHCc/p8vWtY+u3+2zMM56RPjXbIdF
cfTiumBEiywRj2FjH21pv8GdX2r98pWSdBMLvoEB+Yc5PIZeFzwA545dNosMcbC3yRqtkygsgucd
KA+DUFdcJwwY20Hh6yky6Lsn82r26eBHU87YbQxSHp2Loyeno8Svh+lh/wDe9c83MtPrZpMDELXG
yCQvvxniGFVIbXLNEMdzi8XoD48D+Xv0nLhC4fMWq2O7myGItMnnAI8/ZLnwpfGyyxVL8rJKGrD1
vKBns++c7QTX6YTZ421mNVm2kAQXwRlFh61A2U+hU7LQ+MWMX9I5Y3+cd2E/8bEPqjIILqxVJeAV
NHQVk7VRxD5r+Gs/sFAr+TXrFycbvxqyTaZy99MzAKMElaGjMyKumj7TCCDImlKmqJS1B6oRmKFy
br91/PoVjr9pWcMsguL5uuKMEiLJHd8dcAzZ+V0Orsm0AW4LgK9TAxN3L0mAYdRHG08HJBVCtdQb
f3mqRxr9zz8JqTrAQp/6PUS8RwX50BxYU+V7INWCE1bapIKojGpJyidxMiUFMjJsVKUko3sNQ6f4
sJki1BZTnFiW2+WCHwqhM7yCW+c5nQEoqcfHMRDVD1wgMtcnC1o9OkmQnZE7mhTS5eh+KoJQrzw0
o2Ok3HPM8lotTRP+xvVYLtFjabvWfLQdKBvEOBlzlb6FsGh9pfn+BSNEdlTcdMbTjMxNunLyzivl
+pJbY8E0cTSl3kfnfPCKhlaTstaZiXy7ze7oMMk0g0Acyd5gqWIuv8QvOkLPwpmKMUwqLLKdOkwP
cQcWFg+SGt1vR0Qf3VWmlY0WLcawS7kStgvezEQoWKvC84SRRVAxdeAcadLhrWaqngNm0+y1On5f
HvAGNibJXHzCacE2sb0ginzSyJh0wHBSRALVLhoeIrz8YCuN3oVu2LiVNOXuCZeyR9pugO4/wg4M
8zM5TZHlD9hykVA4QwTsMcfNWr0KReIjH4qtCZRhkFOGShlzLwsdvjNQpt3NxUFH+onK/VqKngby
1C7kuG5eQv7wkkfQ/681X2J67ZLrOA8z/8vAWClUCJwlV3kyfTQlHj0IpCyoom+Ze9Bhl875crMt
qI2/uWq0HwXVOMGKILikDngBWrBPid6D9pXCxvrBs6SMegtOa5akm2b2FMZcvAClRS45QASP+RJ1
dn+FBGlG7+kjhSiujQGHzR7h7LzlooowUBe4iFtomQPR5udQmVxmVcoWFdNDvKSbuZjnlOaJ10Bg
bf1bijHzn/ZgOLnz3Gq8U3L87AheVvTakzf44nlGN0kf65tTsx8UIKnw+IkPS9S8VvTKwI4VtEiO
gc12BYgyF7739IIfz3i3HncGa0y5Dvdo6P7nTE5AqVPYe4nejkvzx0zsXRmRfp65G8VF2ozw1DWv
rDWQ26764Nk8aWx8P1K2BMSNphF/PCB4VNhCqEpRo8bc2Sb1IfaCLu4VNW05D3ZSG9+tsAsjHb/1
TLKNs7neW6vTeK9Nlbvey2w2e/bToH/0TAfh1ZLi7EgHB0T0j7IZxlRMxoS6s6ZWP2E97LIDKL6c
jlOR8Kd3um8zMT5zwxRNNY3kU1OKY6J9dZM6+zSbLzLqMlHlC/r4kbuK85g1mGwdqSM8WFb6kWpl
jGLoWwLeLo++z7Fyigxn7S44ZB67oQWPdhe1dbFjFK6Wsn+18BHfvbVRKKtpzMXbmXX9OdLX6Gy+
B//OdaqPnGfm4Zlaix90xtBl4/9HmeqxsnBz3Fczs511gFNJRRFx2qcIELHiAGEW5VjkslFFpFef
zgtSf5qc5VlFVeEG4w7z/fO4inYnDaA+A2istcqesJKbygL0t+/CJja27hdFbfdrDGmR3UUd5djm
WLK5RonQY/PL3AmNHSUqnACERYRYVb34MRhjt0CpZRG50OUl8qnbNws+fvJqXOaupIeqA3blhVgh
CE0YReAx9d9aFsvviZ0qAkmAdLiOXDUIAXjIQZ6TdgnQH1Xx5HdEIINpL1nPNUXmokhXbvbPX27W
Avr1mrBEc20ABkBcS7LqC3BdoZTnW38gUoklxNUmC/4Bf9FFKUtQ2kadT2D7cHZHPMJ3m4WStpds
f1URJ8BtL2sqhMBGUSzIK0e6C+OnL/zH/6mXi2GdLPcbA21SDKYaR9T+RR6WoClwZ+F1iuKsVdv6
WIYmA3ISnuUmTUlnBEPbt4UkG3pDx6i1+mZInWs2K5y235eUy4FvIi82i2yoP0gdf4G/XziY1vSm
pNphwkzoPtSQ7mz9HKfHm21HnkPQZXZnb0OiNPPZEPR4qisX/oU901dtpcVIFiGjs09LdtBdLjpT
CgAWOeLCA46vJ/D+lKQGKwK7gwGUO7WBfiPHSohfmDd3K2qbR31JPjUxTC2rikHh6BNVangD7z3e
amkRQ9IP2LA1oo+hiOV5maZNBUdTl9ka0VOUsegOzFgDsLfpHm8Z16GwxrZF4BWHSRHqRpQTxa94
XSYKBFL6zd/1WhUYtDlxOchonZvnKUjvCLXFYpoDOdJj7uQtbqONbpunycZFVgL4dCNIMx6YOwxT
pKfl4LKov4/CPAr5thvrDZIva+LWNa4loOjx/6vP9VB/D6shWHPz3PZItn9YVESwcenmccJyKlnF
pfwDt8y+J42UERWIwmE737/23zZnwT9HRtIAYytQyQ8LAmg0SDf9Ie3Q2ju75wxJt2NVgPrQ5/xq
jRrjqxz7dSmsxzZ6oEX1boVacanvoW6QJVcUfbM80Sn8+elucr5hf+2qAYRtJoksi6rUCqCfVLe/
NiWoG5JwDo2IErox+aAy3mBAHlmoRXFAzSYb1fd3VwniIsdlBn6WYH1A1ty/QCHTFhevHkwrAn2i
gSDtrReucnPRCwaS1d3fV+b1WUHOTl+kdOjMa6nS+aoYrwrynxuFg6b+PGz4cCnmg/oHdDLyUrrC
JLAp4cU3EJw2yvBz9Puq/nYYUDHZyEQZqgUZfxPtdRkBY2sWOm+uVNCjzr1SEKqouJP7M0rXjnYS
ozDFCZvdxQ95YRL7NbmdnVVv7fg6fOTkDlP3rxZ88HvcazTrHTi6cak38Om76ISblFbIhXFOwd/f
9MRWwNx8NuyUrdmJBz5xFjqRUMLcE4CDiVn+hrxXYArkHeoY/COm4Y+q/KirmN4o9P//RyqxJOo4
l1PWBOLfGC7Hzl687LZQOctJBMDZJujHB6323X7VIkBfTyEs60eGAB+4pQ4YJXzQ5DHnSP5Mwnob
MdddBITrzwxpPI/rxd4bWoxxmWwcOocljpPRX1TQa4Mxsa4l80yizNU7YNOaZF5AOikPMWUFPkBt
/rm61KLHiVL1BcJYoTUMcMyZI47UZjO+BXt1jNoG9SDhms5ZlDGKzlYgnbcD15V/6zBhpu1J0zc4
vP1vOJwEmJhXBf/+I11hwBy8X4hDBIOWeisTYHQ8QcJZbR37FQt4ABu2j47RvRcVqJSA9tGQKvh9
1zGAgg9W2sI+6b2LCA2u6Oa3c3j56KHs/TAMYkZ9n74GhVoqv2rVLeIG66msKn7s1Gxpl7K4zmZY
1+BfSce52ISsx4G6WYiMYDZOdHFsdsOv8aChByAnhYlmfNDfvTNeKMvKVf3bQYfYW2RbGas6hRWx
Dc/koI9ycMpmcT7iQeoNCMilIlHJYPruB4croKapSfGVzHapo5t3xJcYZGyJ9wfkK9PYNGXmnwj4
ZTRh6+ryfhTw3OvJ89j9pJF3Ta9zsjHzJbZoOqPh0/Hyb1W7QBkR/a5WfwfrIb7tgTp7XIt7TDd5
quXhE66tEyXiRxKuM8jrZ66oCywiydjnxJ6spafaPRzn7zMQ1s8EEXtU2EECu99sZL+j4AJ2OwEX
NuyRv1REFguSk1er4xz047j+SnhBYDma0T02QqnKyw09/dVYj+KraRryIH24AN/PjzcmYs5a9wI6
H1VvLkmY2IeyQuRykdLAtXWKr5qc5QNO3jclyyit6JGuxZTh84QzwdYNckROe+lrC+HlpfeLqpBD
KUwzEEtIF1UMhk4Tm84qru9OiMiqe19PmcouId8Il/rUY7SUfl7p+xVY2KWES02sZfKwQt3ERsYb
PV0YFZ8I7d/iu66eWyV0CdO3ExYTZGTezkATgx5Yl8fRX71Eq8PuyyleK+PwhJ/RAhCAZhnr+Vs+
OuPsRDtyHW9KRJku1V86jfSNHg0g1DRSRotCbpcNbxlRxZuaFDwGSEwRHpZ6NIcNw2Rh/N7dUzhY
VIZvNR16TI9+GkJq5MIE8AFkf40OrtpUMB9VOHIybyAOS5nPsMC1zZl0dDckNKidfwoIr/UnnAw2
O0WFPd/D0HR+dLhe8lbsurPrhMgJclK9+F9O8Vk9+IunM/xYx9gLmmcoXCZoKB7K6c+GWWStu1VY
eglGMWARtZWoofH2WKxadbPDGmsFDi8Kn/diCPCUV3mDV0+jXRMa2GeFtysHpYdURhhPlPFcy7UE
087WMkBQGXDYYJTFQqDOzDUjh1JPtzjW0NSMTaEnwE68jZyo0XmNSKuvb+FuEjOE9CXSgOYWnRsV
0tGv8Ykv905LldfbOEBs1DCfH6pciHOm/bq4JYekHf7CnIxzUrgywCmGnrUQhKDw+1UHPCTKftMl
XcbAhNfKWhxf6LXaJ5qnjGMOjAo/GBpJkOPejjUk6CH0Xrp66UflaFWrHvqiI5rRZ863ns0Y06HB
9ENv3AIt4KYrg1mpp16KO9qHWO9Bmh2B3/ZsQopD77hLW7zivOnzgUH2cvEosksaG7owFHT6Jbxl
hsUiTGRQquAvxNxuOAFBFWJcXTkwdgg/F8SURgcUWvprGT7Wh+qksyjsjOZpTvpnd7FQeXsXpunc
LCi8MvWc/8VVVGDHpxVP9XlekWU10YtYTcNWVgwXWwAe0zP9cPfBHuOLe9bIKgUuJc7fxfmUdM96
o6PVkCbkgfMJtfVD+KfhYWxXAKFpMw0mJ9zB/0s77MJxDDlGWG1RGH48PvlmpVBFgWDYb4iX9zQ5
iCyab9UAUqrmyElogp2lMBGLJ1ZqXFt0UBJZr73NgOjGkxJWGfnMhR9BElftfDgwEyhWlVb5F1F2
m/MPvVJheRdUsj1An7G3nG/rm1iYHNPTMfCum86KEa+3p66oI9zhYe2XFKxB4sSjnMiNuDurZKIL
53svkN9Mljlp9KofaD34IbpZxH0FJwFNTfmtIfOhOOxjujRYu8ppaW6FmeP6Arc7EX0qUFn2A7ZS
nlM1WKkHkHxt5gA+rVlL0QUNktvr3jmKfGKKTFKhTd/9B5KAogCI3TUi2HVyrFUYpvUuWzwf8D+1
rmRo+9YiYxzrSUKu7s2FiS0maqyRP0hIR/W/IKkFW03wsvZZ4dBIyx+3KBYZEC4Rr/bEvKfFqOoI
+Yr9XcI4U4FhWnmwh+VCRXApHzJUDhNaPtA+1KoulZJDzy4uzTrNLP7uINBCS1k6HOt3cCSQBuOC
RM8zCstCPdCO1MJHX+b7DLwQB4Z13YRVzeu6WukTn6KaNPln+zoPGr5S4nJwpWiicfj/aDp0/isq
DpNTdwHgd7mF5NdfYAIkX/8Pb1CDkM3sWfODFTDRIFBftHa/4FYkWBKZSYjW0wwjF0qHtf7tNsZu
jC1R9Og7bEfNOlbN57M7iAe0XHOrD2YmlhLWUcLWjdWdeBtVl2n5j0NJVbFTbVapuUDi2E4P0NWk
imQoqR9GIjyDPGr0YDjYA2qcCms+nB0fBJ59i91KRh8eKJhN+dPtOHTMuyHf+z/KHkBvgxawdSkb
7caZmkpV/62D18e0pBj5eQxdQyhVB97Gh3tkctpzfB/heDhDcjYOxnwqICGo778D9VBXCI+oRtz5
GoE2lqkbSrQyyaQ7Iz1+1NW3xg/r6MspUArtO576VdINhBkW5baS2OXI7uEJEvUW3qM104KNMHNh
xiDGbeGx2sO+jDywCQcOftWwsHSwAlNufn37sM+DL6RUY6tNL/Ulgkkq1UKiiMFqFFegeV8SpOZD
ZnRBsmx5c+WQ6bbJ4w1IHwi4E4jVIV6qosi9qUgyLOaHBKBiv4OECkd+sDwGLNrReHUo3O0qq86s
y83WR9WLyBNBp4aTVE2LVrhmJJ3eeOmJ/rZ7sESl7awrD94IIuec0UrSqkgfCS6VKZpOffO53TJk
bRw7i4W/95+pFch2nX4UT/EYKnqTUDQa88E2tWA41c9Ht5efKaRieDh9Wz+eaCU4uFU14q0YoCOx
Q8LT6mVl+zHEB7gcKUqFaC1sPX7miRtuMpWKPIYMsuT4SZMMNLfDfBL3QdJZOzzvGg6lCV1zNbSG
f6zdL6onbX0k75kUu8xXS4Drv5UBJ/fhCCyawlkjpHN9pL3VdM/YvMpxI40z6rbzbk/AQkxgGe2d
yklw+Dq+12JD2X/kBPF99hLXTZNKRHtdh6QwIIBpKX5KXeWmYtxkWgV2ld7ksfBR3mNr5kn4Wsn6
EjyTZbGdSDH1cN2kIe/nt/0+gMhNkIMWqY1qa8Xfq/XMoAptz1KnziCv/9v5NhSBxSBS94ipCjkR
aIppFs1Z8w//MjDxie3K5W/1xsr50X5YlTRIffoq8F3TBfVS47AyRlA2PXCJaF9U4aEpXvS61SMi
5P1ECNW2/iwud1Zs05jJO2fWc8IEa5RI7uW/ccVwsDGx64JaldBZqFyu8pjMZCG2tZkIYeBs3l+g
QghxbjHXy1JlH8Ln4jJqb0kwegq53w/7Ot0J1oe2Zv2wbVLu/txfz5JNWIGA3DcDLa4ZXp7fsgKk
YaF/CN/TQvAnBAzi5RYWTTYOmUSbU/IxxsEB8LZhg8E/Jw4uFpcB+8s2jADLcpOjeNfSlgYUbkzA
ugL3HMAb2Wubf7EXA7YkzYXzwld0qoOHcPT/cMKpg1vaIvjH/or95Dp+O/oa7E+Pcr6yhmcI/vkQ
06iVkecpftU2EnYflLOnXp9fOIdCNG+Pe9Gl7pGtWPXAyWxxWMDbammB/JSpMmDOjiIuxE6RLoAN
DJ/p5daVFKE0dX+Tdxm75Tf5JtWlkUtl53+IibQhJpWpkLhzLurpq+TDxhE8iW/vwnxVWcqt6zFQ
ImpSxDT8r6bF5PFNU0f9Ub96LSDW0AT/rEJQqH+2i4v1/VXBYjbxDcYVLHXJo+zaQtya+BS0ZTkJ
56yPJttvjMBNb4YeOfon37QrfPYtJWKhf6zieG2UR/7fUep41lVZhjc09ZlQ+RQO1Qnh++z8AkG+
lEtpsoHmoajbhA/D9HxsxwvEqM1ZCzRHjo/WXDhdEhhfgiS7vnjrQUDmf7mlr0gOIxdoqayDZW7p
MzpuWtPyWokkKlPDd59hW2BfVzKRvC03xkfPW+m9O7pcQp84Py6wLbLJ8jYvzFzEj2VBXG7TqAdO
2H/ZQpyhU933+LMXc0FVe3Enxddjmt4FnxMHTqVcdIzHXheJzJDwqfl0OcEV85k3WWneWteI38Fh
qyT44YqeEWxBIkApetfC2zSbfsQa0Wvr/tOY3sfq1KrcsX/OFjly+txoGbBHgTfVLzVBEhJ3o6o+
8Ro+kX3DXnsaiH9W1dPXcLsMxj3X74pdGFsAKTQm59E4Q6YxQiN47SKyD24WPO2w5RG0qJuyVpag
wyC0fCaJGb5x+wA+0SPGu7c7fahPk0kaU549RjT08Ifd9mTIcZWgO7Ghs1d9T4Jy8VobHT2AO9gn
/WGT8JIOqI6p+kBKMUDnVBUFYg5uGY5rm4BLOTXCl2JEQT4nYnazdGxaeF3lw1VqrD4He8sgjNts
p2xT3BNDYfWIzX2hADx1DCzqnm6IuJmH8pKWwFLECeAlMobK3YM1uf7xxj2FsCEc1zqQ672p2WYI
Tc0YIrRpZIsmjigLiSuUIsPjK793Ydj3YAKoZaCbStkQvnP77GWBurqICpHYE+9putiZ7+m7VohE
vXxDrG3aDwjCxivt+w/avUbrVL4Sv3dPUmLPCtsevwJfoEAuck1sperZCk7pqo2Ej/3tIE++eJ8L
LnWzbFR62VQIeu/d3np5n9ADdXto+0uShiZr6VJ7YuhloD3pzru31862OyG0uHGLpOut26NPAWHi
z6VaWFHDT8fL33D6XBLjdbnXjcb96/IirXEC174diwDMyYhDcWL3dFdKpUWPUOjKq7mh4wbLy6jQ
fvRaJbbVyi3jDqMfpnAvnV3XVdy7HtDbP5ijeZxSOY664C2vpN/6br0rMS2chHAMq6vjSyuNRsJ4
9bpIMwSL1+JdpKCJKs5KNvMtHSXYwySVF2pCCw+ru5MBeCXFQ83sN6P6IQYhfm/uZAYujwBnOEJX
YFk/gF4nuSVr6Ds/pFNCO/O1SwUOdZYOEs84oZBsIzoQIDbSVb4Y+rbQvyvKZb9A5M8fc/Y7n5AR
gY1ZwMX+4bqJFA7BUKzkSNiJq8NTCmp1Ok3LioB1GaonFnq+gB0M9F/jkCJ9DOEhT8tBn+KIbRDn
kWvgg13p+K5SlDBg+zb+lxYvG2gHu+yZt9Yl3IcNMvL3K0yXH0BmpO2Atr/cjVuRVeKpv9dz16OH
aLKWM3POlhYTRgLkd2hT/Qm/3tjP8xd7afUduo9st4JUAyZFskyI/ZyVbhM90mqC7Qr+5x+T6jNc
d27G+lZA+IXSF69GVJWAed30youvw2GLmmeouxJWxisicDeZ/hyLYCSw4hFUOsxXmmOyqGJYhOzr
efl2f6Fe0rlpqICEbmxoSfcRumCdDK/XVdJ+c21BnVbOi4heuj0/z2wn0aDIMrQ20SJa8oTlKCnu
JaM4rYIlMqb12idWZ+FxuzYpcQVtXDWzmCx4ueQstrYhoyQ/dBPFPn2cPgh7npojhtgUW+Ywid69
bDzcmbtvkq8LkiQmvU9QsYsqEhb3ckJvA1fzXZBh7GFx1y2Lz0xLMHfMvmc6p3XXA4upJt9rYkNM
I6q2qD7liiurOVcNAPLxiiuArRICVIvoXZ0n2Z0Vx1HHcze3KRouNAQi8rTNqD3F3GCNCjFzJDOi
wQmBjyXVSbZZDESA5RueCoM9F4U6VcaaBiGzo2zw7QOvcy0p7cqvWQaBJtYX4jxWrL2vqIMi5CM4
xv+bPJiKFMGTGKGjTJV51uB0Vyb29s15j05QpGgV64kFarr5NiLXw2J+XThWf6ZqbFXizb1XsK9z
eLEt+bj/ZogAUIDbov4lwgR0UJ5DF9xMbzszzIDcDhcfqqBAa1Km81/8vrxDSqOpQU6WwrJiwQxr
i03Q1tQDUxd5TEHASHlCtk+BWB2KJwXAhQCNU5Np5GePpaqFJICBJ3AtD0phaHUp7w9JcQ8s6sfr
2vxQDJctmoGJ+kq9xMdFK3HV+QnoaeBKncFOTpw46UFMSixfArq8wtfKwv1ID9qwjtC3FIjxZqlU
RT6pvi5CMkvzqRAgOQ1Px4GfgAQlOYJxdMSsdQYkQjUTskD+65uKrI4OVeVKPOHlEWFQ0+HdQP+5
AWkmgBDGcODhoegQqHNRz2aSzIhukWG/1NBl5QGYlt5Hreff6EsswWgONw9hl34dEafWNTGBxDFU
i/ZlQuUgdKY07o/KBZ9LUwCPyNTB+VOoy0tJFcu10I/AoPq23sUaU6SUMzSuZY6EwSZrrWnnlQoQ
i1+/bzdXirg/8SwxIVp0ZsykEDBqgc/vfnKxoyNv4ytv2VX8O6QMU9wnhf38wwHR4JST3+Q7mHyX
Z6WjLl4OyX7JDXdSAwY0CxfCUS5cpPaZiljwMoanGZ7P0sXq/Val1t0oe80z0ZwVIlHZsRJrsv9E
8T2DuevuCbbGyHiHd4bJ3J8LLdBBfPtRK+pKIBj84N2XsvlO2CJRHG7pV4gObnIQ+kkEu1iUtlsy
wLOf3kpxAxoEngzZKIZBDXSYxGA05fvkScJEj1OhHotB7g89ynNyzE5w4UXSHMp4KR/8PEntFkiD
rihgLcvacdGmVAmcjhuvYmgZItv/IzzyaKGC/CyFZp6oevuKWM/G8XQjM8/WtgKm26gEJjGUgYXf
JuLGuBv6CKACfutDE55KmJWqus1BJ6Aimy/LeA5k5SSCtDREiKsDlCKE2tq+IC0AbD5GtlUREf5C
qJgmX2yg7lA7rQHab5ND4oFePxRsLWJMmZk+VrosunY6urKmjuEKOHYZbuMgosrAMlzSrVelei1v
hQIQ2Evyrg7qc9dI8/wdVmqMu4ifwvhAWRNdBXOEgflwM5MiuXjyU4Repwn8XDIOzKye+U10yPZd
+Xz43WgVbjMaWzp9wOgguIu8JflxxYLu6fyk0UlsGgiXnlYEHT+my44WJ9xeGarUl9JeP23KYJFo
wCLDE2z9O5yAeLwi4rvBq5lMO9uW2KQ0YvNdmzEQ/VLS9wn09iY7RMf1M/uKNkqVfEiQU//8huEK
skXRSelMBifkCO2i91kc4a7QKELAVGsJ37ZDwphCpd8y22yPbMEkzPGqBoDJVo2DePCCkxRC6BUl
KuCW2t73xiaP+dGNurl11q4uEf9xQzz3QFtZw21dJoiN59wjtWvU8zHXCqtmBgLae9kSh2HoU7Z2
WqG2u/aUTCkndRasx9Gwn4nLvskcwJeKUiW8RtZ6rak2DmHmF6K/JG5aXNdBOMjPxr3JQwoSQiPa
GxqzvCxhfIgdKD3mohfZIr/toDPOriE1IKV6gkEiCZFL/LtPvdErxkUi7SKsN/Vuvp5GEG7ISIvr
GW4KLtUwvHbyWvhNjHYknyaFFVlhBS6jvwTkp63MpjAciRUjYG/dupuZjh2vU5YXKfW6/h7z5PN1
1QNaWHPJrp6X2HzmjHNKn341lXG/b3ZBDtfVg1QyisWSwqTX9VfE8XmQKaZhXGe37awc0MbjlTJP
xFSDAbHc6sSmp6Whs3BsBFu6ACliDc2gpEjMuKjlhwOZbJFBg4YUBW/6k6P1rMWUwDKw98LH1Vzl
oDwLmTtMIDQNtwQhGRwKlOksfRa5iXcma8dRmIGkiKq7IXy43rgwA2GIEF75IY4npCNlvKIiy9c9
rtK1qwT9f/7bFxZSKX5B68YzOwkoROAfNCnH5taY8s8GV1ZEC9TrbSFwuKG1TtLwTAEBDB6VhL5b
oKsUekOlSEDbSERidfJZJsjxiUf5t6swd27shTGRJ8G0qPcDB8+0AinJTJqUsV5Gb3LP+P7Pp7Y5
sR4BJcDqsaR0vc47tzanwMSTScHwkOdnYoJ9f6nZN1NfLuHbX/cDjgswlr5i9DBfBxmhWZjq6e7W
vNekM6kFdXFp/tdS5Lx88dGfV8fj2yayNgIlWE9fU45LFROe9Lc11Ppiy3+FuEr/8OUMYKqWC1Nm
MwrC1GZ85/6lKSrWZGLw1J1QC0bVoEjsXJDAaj9TLSp4rW406q9Gdmeqrmg4YBFhH+52nhPf925B
DQIWH7uzwl1njy4Dxy4bd+wpi7pXxu+qw3p7ICOkUw3QgHtKISwwdZjy0fTWW0zz6zpVle84GOvp
hM4ZTPkXPn4e392pS/a7/IZJox+rpL0aCKtrOB0aLdPb4uCS3B83Im1vbmBkOw8qZ5z1cWxW85ze
O4LHg3ku6JVekDFDgB9LhQS7JEzLTaq2fTv4yKoYB8GAaDZYTUdXiB3CKqgrI+vX7aXesz2FMft4
zZzekrrNRW9g/Qo7+X/IWA/HuzsQqFn6smwwx6rY1j+/T/pC+eQ6y9o791k5GaV6Dq571zlCLLKh
jbSkrJgiSMjfBPsIX+SlWICQM++9QRJAOwGlSFuYjxY69gJRtg1npew5zZHX/JQh1VrNZEtKCkTr
jtWuIHZr1mvTDePQflMEM07nlSYlTn5Vim4BjOdDBdDsV+hVHGEeJ2aWhnY1PC2UExhc+bFkTTwd
GrwRpvIM/TmRiEjmRwqmlML90f7SKoCpR/cmVvoIOzq3SxTgjKky1ui2oWd1DYWYajnTLzijEbPj
8TZv8X7nBqyl5kW4kCs6hZBgI1eYypnuM5MGfZZtdJ56+zq0BYu1s0iPU08Hsv3WMTeCi9Y+APcH
2FeYfp6TpStylf+4DyHpCenrD57vShtk7Eflw2Haq7jT4MU9vDGYFTgmKamrPqWmcv8bDnZVuRjd
kMrCHp4/PGLkudYr32A1vY6tj3PWxhKTtFaDZgjxEyicSG13+4KB5gEgMi+S8KEM75cO2Q+gQWTM
g2Gkg29S03AvGDxAo4dRkP0B2+Y+X9ZC23tSBpgMuqCtnn6GU5pqV3K7Ak6WO+/nZNFqKmrhQvE+
kcvNz6makk4oSmuJ1/OmBjDUjLXfDlcpW+5WQr1UJ0c06BAWIl0Z8Xy/I9PVf5sW6gKPa2uLMB3x
nkUKWXKI6zoZ711AlaFtK/n4Rw8+xUxyedZTaU+nOO9+6h/KBv94gxaxYVVwNO2UFBrYAoNSIG1F
gZxCivelTKHgrx+UMZvrgpu2InCYENsuFm7TBWqtTn7kNtswXDHesWym64rGICgMmsjTyT1pf/w2
CFM3Ieufn2RjGXWF+xTBVMjZFPfbX129KyT8STYn1U/BZ431/GDIfdn/eE4901Wjqz1hoDXk1TTr
j1SwE9Ct7L3C000bZPLMIvLGb+rrxuazWZQhbCiw7CABhyDk84gFX6Oq/M0RjNkkASdw8d1aypFM
LK/GmkrdZiMXguiNMn0DDylYNLmqisc/oQdIefTWDeScbbqXXeS+IcW4/PqLdlRt1BQVEUKmEymP
RjCgYsl/p2wY9ds0IwwNJdpb/okNARFzq1bUvffCo9fPr/y+jbQmcNdBpl1Ps+zUJ6821LJnRiql
6/tI67hE0qO5Y0jJKaH2fRoPgwHdSyr0NDI7sCfxSaDAdKofirrqLEAKjD7xooUOOqBepoQMYEGG
zqxE1SM1jtXhpqd2dt28hZ4X2awTCIhwwWSx49v++MhFtluRbEvdNrtTxY+fpLvgx5D++pda933t
NqKcYPA5Ho8EBl9imuwVDDrIP893fDt1OKgCiSGo7eQM2IfYt6XNWXJcoItAxbV/EQpCsrFtLmU1
jkq/8IdSMjCXy8kPo/mZUO3a/5xcZXKGtJYrzhxyAFPIgSw2E2CK0ep4t0n0BF7QUyA5baEydU5u
uXwphoJ9xAjD48xDJkAPbWe9AL6zZ0DB+dPGJn7nuTprsg/jW6s9Q9PZeGNKxksE+zu2k/K0gvi7
CWekwzD6cHCKYXe9keus5zcl0W0Tbi8srA1N+g6yRfKKFXTee40M9wnmraCtS5F3U3f0h2aK7IFM
u0DwSb2nllvQi7xAzUIZzHOs6ghhzDtzDgyvhFvXD53P3OrtnHcONGEYwHBM3XBsaZ5abM22ZHkR
lZvgT6oQHk6lF3pRHPSyqObRM1Z3mj+6tdqVRngJwDBdm+JzpnL483J+UK/j0beaPsDvrY0EYj7x
baKPeVkT48ooOGyVDOKB8P9Nlfek6pC7luge/petRAK1kT3cpTKjKmAT2iNbgGtFTMKKTYN5ccdR
OKeNoOsM85Ip024h8pMrDdNsA1jIOEBqoTn/TMhjYg327uBBhFXd8Tm4Ptbwslbg/EOhe5mPbgMB
+nYQAiDnYNQcBxmfa29UjIawbsKm4CAvDK99n4d0hnGQBCqDWrHquluKchtytDSQnuBKNbllvlRj
fyUjeBD/reMj6vJ2xck1MMn8xmXTPVZWIH56E3S4FtPqNhGSH/vsWoYT2rZzM2fK7wXnFC0XTFwi
0C/qaWCrdFCa2g9lESYoVFpw+2HqaLfJoLsIcbHJZ8dUmRujYuP4HLcyvkO0JQrcSiDYA2zZMQLR
qXyCxvvb7C2cUE98cg4lUC1VrOYxYsf7ifPAAf7/3+YZxAjxqQa11eQFt0Ml6ezvVgmqln2/6VUW
6d7vuucgAXJxtLQ09hDeh8fUGU9485kNAyRys4tDgrsLiyRT3pozJCLURSGW0NkpkD6HStYhrmip
sg66EnSrzd3xdfaKzaEXoId2FOitx+DmYJd1sX9hMQuuZ1Ai3jCa2FEXpycJNZshw/s12eS7JMc6
YyyWwY2JjwBaxAtqZ9iiSh7bq0XQmXDov+7xUBI+fXFFvr1JZqAEE7dXH1qw3rHBDIe1MiedFGp7
ikzvfTFb+oqvwzfqz4cm189zCZjkTZpOaGK0l0hAOhG9shw/4aVssZy6T5Lku5TjD4Mr2cgWF99X
bgCVUks2uknCS5EqP0Wda5MFEkZNSf4ViAlbP1nKZHwo3AI5qn2dHtBS1X8g7ZI1Y+g6u3QNethS
jkTDaRsdC5b1f9dDJFurM0B1TGCcZeY9jSlZ0H4i+3fNRwzxs989oTrVusgOsrRMHVt9Mg0iOiTQ
bArt2TIhiqgLrfQMF6BfZYwnV1YF3Fq37UCqogpRM93+95ZxnNQ+j17DOZka5PGIsWQo5zvWGDnP
JC7X4fTlR+cqC94dWpyK2G9AUY+M8bHnyPcRxJQeutc1y5ZxQ/3XaMRNtIYdjuEmfzMTGFtjKvbg
lhBBJIH1xLoy173wajg8iOomhDj+wRenIkOAPgEoIpSpxbtlQ+sBtM9x3omQm49Gkeg7T9wUm6vL
Q8EQHHDZ3q3xgzjGafvmPhDnYKCLDahfazbxhEHdZRbNAxO5Gh7s0wjCux8006JeU4dmwFYV2VYG
LUV5bqhg6oFz0Wm4efCB64xZrpkAx2vMZC/ZMQvnE8ab+E+sP5bH8hMGECScgkYGmkLj1w1otdgq
ish+rR/aGjRTLPi8/ldZ/PM6X2ZjKpvKTCSt/MQLA+0xLrX6buZS7eZRYWwtY5uo9UGf0p85IpEZ
RBfG2Y3nvDVRGv2PYCJTKWnfPwQatUAI7x3P+/4SUehSNIYk11KXoTjUVQVXWW7Q8K5bFtckzocq
JxPWOSRGtc791xcIIK5F9rXQJZ1aDnmhHnaAl5PCka4JmfX6/pnurtwXIwTQW7MEhqkFIP829Mne
QJwwfD3YwCuf7UsxO9ioJaCKCP/vqyykqoxTCbhpXOgHmsXLjj7VQ4gYZ5ZZy3rzwifKSe2tyP+u
935M2LMXhAdolPqYiIHu/3XBkT3SsLuyMgrxPkDF6glE0U0qfjGAr9aB+qz43cXs2YI3UIGa4j/E
Lfgm/hlHFXfkfazU3qQ/7c3PRug9iSEO2aB0e0SIEfpc7MNWKDbWlHNNO8B7rc1st3LtDfKqYoYP
/Xac8mBIfrK9bABaEa4CexVdY9B8P9K5bcP0PBJ2qDy4ygio9sU/mMnA78qiOn8ypyfMFGi0/qG8
Mf/k8wEGUA8n1SAKtmh2XyD9n49vBNpuuWJ4cSYK86kkF67d9WeSC/6IOcI9o2sCa9XF2reQ9GQT
vv8fLFXM+WJ1pphjQlTWturodzvnLS205jiILhjdAUDCk+oKJMp1gMjpDntvv3hvhCuuqh287os3
lFYawmC9xnCupHHVmL47iVCvE1o8CncnJSQE0KCabgbB8aM92WYskh/craAB1aAM9ozCud11AB1P
yK86wGzqRk0pR9USBLVX5fAowtBB365tlnoy93gZLefiNDsX8NU0V0QD9dDfbk9JZn3q2cXocWKF
QAoPP+mtdjMQG+3LmEC2iESaJNQJOXfC3NDnZ9Ys/4RKAllha5/dqRCLitDuEFK79KqIEqd6LmuL
lztIdKF8seGEi8HEADKQLpc8l6b3oTTsctYHf/XHj+rJ7mmkQ7QuLylWT6sL15f3jinZtBZ3Z4rV
NabYgnEupC0Afsw/NlNex5PmDLj28w04F/zXm2Xuo15uadZu2axEdP/IhWJ23qS2Z7vnDLVTyHL6
HMzqPqeS9b6zoOO4C1Ht/VgF+G6aLKJUANp0IgvDr8nIyCXt9xuaZit63TVrw+FN/+cItnq/CCHs
c2DEwEteI2d9rpH9QeuTuRdZGX3UXoPFl6UjOgBRzGynT3EtJ9nkgHMaKJV932SiuY5pn8KMSVo1
y1YJFNoSCtHIqC+rwf9OGUcR8yJ3eTNtRFRkRooIRTpXZp9mYq86y435tkNuBFbDXBBk7f4CW3jU
V/w8FuqhmjMohMn8P+Q1R4c8GseQSr1GAC87An499S9jMufoR5O1cpa7OJX3j/++++la5SFwpuXS
+YN06Y3XSFlE+CubfaxAddOsboQQs0ouCQjQD4Wh+BOhh/wo68tFD7ftLh6OucLdAjsKm88iFHGF
P8OJniEZArIj+KKL0s/zp9odW/P4Xf+me4wM9N/2vyXOjhNbdvngJcIOhz2WhCo29sgig9YIutzN
qV+lC/rYAO96S0oTybVMkzxT+xiS9FWO4EvLK4myknbJ3CQ+fV7eaIYZ2JbyRwcV5AIOQVpdIPsC
6lA6Ywqgcn/Y9oU9pbC39GTF/BtYe3I66bCqJ81OQtWSHQ9PKT4wuTK14GAtPL1HD7o1NthDlL8Z
7Oi5ocQEPKgOPvrXoPGZEUT6X7KPwGVSLDLX4Lh5ta1m/KKAG597Q8Wegezt0fKlXRfXmbq2rbHV
shZ3DoXtkF/GQZpw43VYxKeitD/w2ggkmz4LC6QU3g/EqoKwlFkJnP2YhxxNiQpPIPyfYZKlCMys
Y6hUNY3Dz79Lr8hvphBBxITcumyTClQJOpTV+a+nv6Y4iYNxElGfD6ouySOjmAF233eHOpAQtMlG
wpM698RqGnTHM7RFoY04QLz6slINC7K3QscHHlKw5ja0SLlMTXbWWBL5XyZOuPUrrOeGNtkpAZkd
7Z96aHIzW0Y4ptuUYTGCyxgRBXKnKqxKtIK9Yg3JBTuEqlylG0XOGpI6I/rEtXiCItFenIJn2xdb
hVVE10gNYA7YPumN5kBXFUZBiyHa6F+B5VR0Zfz5i2jSOhwFCrvij2iumRXSiS7XzjyjUNDNg7ot
iCxFZZrH0FOgMpUGtJwRW/XqztV6uF9jlIL0oUeofErLKtA8CKiSJU14Ze5XQUygoSVDRmjZP03c
A9ftlHMWfsdJRGJI9ptjHBh1iccnBNf0sdm3u16DRnh+LX7DoEzYIJPSpogGQqjl1FI182xhEcl6
MQOiCw5ehpSBndQs6ghAacKwnRRopO1aG3iLhyQ80ZxVLOI+pU2MgFcmzkX9ko0FlMEEajtcWknh
sCTscEtp6hzTawGOgzoPjba+pVR2TcpJlJkSUL1p+ANHOxfG4Fd7ArZutxISaE9wdcKsfMJs8p8D
IkH9XK+Frc2NOHLNfiY/ZfAZrQMHIUigNukf8TMglxHfdwtKlnUvqwCu0ZGvgSEN46eADjTYNUVt
4faIvk4qvSxw0KKQNxRXOJUu47xzu2UM1lexkE3WzaPviyUuTtmZLlqXEhqNx1whua0eft9CKagU
rijIpRoWBJL4tp22I9sGI/A+20EsiJ1PtpGNSdyNobQTWviKftyLjWu9crR1T462FwEnt3r5iGAH
PrxWOltVJyR5u+mTAlWrgFa/dmc1tjknkqiiFzFfmGFu17RIken5FvJtGW/TX0ywLq28Cc7N8635
Bx+uEw/ib9+ogyD1r9HZ15vEIHwW+ghVOW9NY/gj3+WX00rZ2mBwbrF5yiEiXrPtvzsS2MiUYRRA
kldzTYl7jMtc5V7yt+Gv3jYEX37viFJXwSuE4qLI8EcZUJ1WhUOFN4mlxynY87jlxr+SjN+HsUFl
6pUeF6efuFdmxE9ovNpySRo74kWatplDCW7U0dwNSgOn5SoDSecWwVBXA/ijyiryREZE6f6v+uN3
T7K58sm/07LMMHlkUooTg1lPjHLll9mzB2In7ZFK3WO/AXPqP96oXJMV/Lwew165GVwaEPuCrds9
7hf9PqbJOjh1y7ubJVZLRobM6zJqr4EniGSj5539Y0PPyGDObVm8XfrHVfEtri1T9bWFJrNjEoPO
ZdnStAR3S81khibtrBGUFFZild/ifKSn+QqQBQkrR2kupHw234oSigy540o0gi172jV0sWYVxfkL
Xkp2tNrarKFCiIiOCB+JOatHqsqybejYnUjQyNhDCvgA7GVEgkFyis4rKblo3lAb4NIXG1s5kak0
7u8lBldNXqXQzMGQHHarxA8Jku++5v3MM8hIyw0zxQzY5P9BkBRyg4FEGg9iATxv5uekQ2L+uT5P
t29a31SMRpUeujLGtQqVnX83KMVSwsu+r4UgGt3xpaU0sF7jjwodkuJZd/dXk09ZLUIP+wr8rKxH
wzpzxRFRw4pvkmadSqKer/uviBN3+mrpQKVbQNtj/1bkuX5lIR8dLcMs9U18iTYRriyzFvoPLgYO
UreyNMMicGcXSQCs5CvAF9d2TNu7BB42hD3y3YCdWY7QLXwAsPUMtm7IRKEbuNUza5spu6F9uV9+
azDlT0wj/t5z28Zx4j73m7twSSJ/hy4tQ8Zv9CjeOXU7uEZ8wLUsIXxw6DPUac6PbeIt5vf2j0Yi
vHnOb8pz9IVjZMIGKLt+ytDJ5j20nU0LTRYpCqZ0yE3haqeZqnHt9Qs8G++7cWqdSzWNk0JwjtO5
VNGJYkKwijWstRqrcKR9ydyMmeZC5Lrw+u2DGfGWB20LMnnzD5wwVzVbhg3JgbMRVZzlo1rzqpMP
ivORncAIZf2rNvMhm0wG+mAMoP0hbNntLkhhaWlLp2bi74zJxWbx+5lIGwTNEEICJwNrxJbBjqU6
Iqiv2izUHIHloMGWKM63gnFDABec5BeXemk1sCOjkQLDrsUWSGFx7LOV6jdmVFSsatSbahVAjTA+
ieLIVAOn0bh+FAcL5sVQvLTRhgUrIdyery2Sw1N53TcIyFZQkaYW07SPYZ6GELy/83tA+WRWB8S6
z5TUem2pSTngj8b7dA1sHTKOsGHsmQ3L45Y32BGEk/eKyAmCSsEQIGAZIytaiofaOHZQrODMfbUX
P+8EcKwCe2aUdCIL15fIOI8vl7zsLLojrlNKc+hhB/Fc/WFt6hsetlX0JgIiR6kVfz1dtZxP822J
+brlpybhPMGopi1NaV36KGF0MNW1KCVysUFf5pCscQJGvTEItCkpPe+iAYLfk2UBGaMCdXhaY9ZX
jwRMWOM2igBphE52bAdwOAMRumsnU3kIBEhZ1h7w3oiWZ845u0daUyuTHlyG6A3kUcTok26IbfAt
7u2proTPwDvJtGln5bLnt+MC3G4ntodIxv2lOu1FJvyXnYubIcSTzPmjp39qo37Zep0dqObfPY3t
y0kqVB2RFmSEt4RcVnxicYwiXM5KnmyCm4ANAIlTiYXLCp8JqEEC4Az5jNJ1gESZQjdWOWjyEbxH
Igi3t8NX1RZqLCsNj7YhaBhfiHfedfIvzds7W4+WkwVlVeviPgf6gkolRqhZOZvOJE93j7joOnuR
kkfx5FC5SvzcbzThwK96SC5qUNhobzUMUP1TvX6MA/3Tc7BwViluN4mZmWiuNDKVeIEC4zz1AZSA
1ruFRQ+yQt1FqITWtzwX9rn0dZGZL77H9/vO1Vm5iXDqbsQV3t6p1zNq3IMwzVfoZLCxzf4a5m6Y
TsMyHmiqWfrFVbupD1PQKFnT35IXvmmEUJ8WSwk7e7yXEKs9hfISqtMP9zQacqT2Kp0t0d16YhBa
lpZ+3/SHT/tqzr+X/9EqGaSufvOe0CJ0Y1UgwiMYUYlpmyCt1d88z2CAkhh+HeiKXDOC8/Sz9mvT
xTG072GVJ7pvtMWVCV2c3ePhu4yhN+WB2drySS+Vyr6j4T9YIHe92iF+cJU91fePnI18/yvGPuir
w/935rGn9SRt5zhRpRz2/R60P8cvn0AsPCUVWpSiVe/0j96Efxt+3HOzW0bcz11icC9cicSeO8Og
vnclaBH+Qi1355BPxKBiy9zIE1CF1Q2JrfYSPQOU2fScxhnhq8Lp2Qe4RXHRHtMFZOU02KD4shef
RSmDSy6OW1lcIWF9Pm7J1RLf1Nac5hiiAAKC2MPrz0oI+p/q5XdFLrj2aWUoTtebp65Mdnv+/Axa
YhiKrKbzRDi93LqQx6XD8i5z5+PS9zjOKSK/ioMSV7DiPVJgbXrOM4wpGG1Y+yixgs4B6TFMWXVW
ZdqnI5ArkQh0FQz2xsxcLO3x/H0lcmRnYJRhdHAGDpNB8crbW+rPr9hGZXprED2AeHc09JQHLMu5
zExbbrKK7SsyeCfUbKzqb+TnyfZHOr7/+3jOdM5TNg/JH9wrhtXCTgT3mmaszgKyXFG+DbRjGO0H
Xgifz4HmtNBKUWLRGngII1gda0AsnZw7/rtJCyWUX9d8bAMy6W89dP/S6p2V7REgU1a09fxnIboR
ZYhH2b6R+6eM0YI1TRrtmoCU5+YhSEjiA6m1dpOg/3XsFdghaGMK5Zckz2ACL6MkYdzCBI3UH+GA
ObpOKR6oN6pEF83pVdUJ2ud3hy+VrdA5kOCPZLRXlA6N9D7YJGSmgvgdCBeQ2hVOEHKiwWkbc0uL
tYTkbohKbYEgShbbm3i9jQVgc6x8aqcd6IMxE1bLCJyyelYhgYI/zHEjWYDuJHdcefOKazhliynD
EhhNYVZYztWmd0oydV6w8g6BnaZdjvg5rAC0Sn4HfRM3Wjg+jLnoFZu5iGQMN8WdUv/r4zP3ahex
PzyGckmu10wE1XttoF4Zb98mtgAUZEQtxVhgwd6oxAdFiVpV9TPvxKbaLgnGCUNwJL8PlClvwEkH
4DKQ2JwFSwtYLrAnXBShKdmNMK7CpCfBqncIjSfz8fiwihMfq3h7tHZf4/6ApyDC5Mrunz4HxURP
o5xYQPx5c0PQJ8s8idoNRtjMAHIbnyZvh2rp90CxJU4OQ1t36W2wfgeVsCJUAl8rxUjSI/ju2XCz
DLtRpD0JsFBp+/0OVW2MTSgJ9KXuQHTdI0TOJWvxgiIZPnk/Wg2Np4iaDYKcqYL4IqX7mhJPKiBH
rEF8OEQ0hLFQQ1cNIfslQyuvkrlfGDnZZM4ltaHqKmRyH/+wIbaDWfYIIQt3+uL71W+PZ9XUtVrp
tPieXXP+UkJEJoKG5cCwqYoLcPE3kGem4f2zUXpGW+r6YyaF9FKsmya+hWWjgz7sDjRIRhNxhkKR
l09xy1Y28ZTgK7qbjVJXjeHkgOEysBN/ca1EDUdSQHR7KAxPXOC7MDClw8gE1E+b2yw71Q/DlA2w
G388+IfoI+j0POBLe/nHKJAUmYvtEtiP9dbyZ/8Aes5BxErQ+k8UijYrcQ5lHaKE/pYuN0lqqVRz
NvIWviyQXz0CFJlo7crX3PJybLkDg77JnzPZSOLVlV1sekx0FOGhucmEVFbrwsZ8nIz8OH+jcjss
l5vyTqDZ7+1wIkdg/kSgI3967qw/7ftf0VMKjDQXmwhzvw1bG+GcBN6kTRycTpQM1JYiYu2Ea/Aa
wHRA9hF9mp170SWAgrCgSMZ/ycKf7CBu2YIKGOQqKthFaSnucjAnMU/oKXosZb57H5IT4t25KZGV
/sm2SE2SraLFPC9MScdDuD5UVbjoRMWGN8vdK44VrwMqHjEfOHK1ee+fgTDzbjexmx++REFoGH1p
Gwvl6O5f0a9IiU1tZF5abES4Jy3Kircxde2GAjb25MRxG8M6AIn1CUNMtHQHj9+QNg2QDHNV9/Ib
DT3y1cl3npigZl/LBdMoZ9GL5MCnBZHBF/Tnw6n8ROo7tFJBYuZMS7h8kkrATCwBK2IQzuJ3ugPl
yeBL7OL+5pKyRhme9nCcgNcPpSRYuBvqDcb1+xOjBZmRtVsPMb+eYFIon6AnefU/yOx0IltlG0+3
JUWByMZeemh8soXu3Q115dWdwk85m+w2TWyZ70WI8HlDcZhbDLFTQ/CpVHAvPPvJk4XtGL4jSMJG
RLvNqu+CtyHIKjjHDKvfEdxKYBzmD3z4Be9bA23pxrR8BemggAfv3SwxBUGoWmUnaIMAUj8HRd2/
Go/kkWPodXvdOol+sLC0xugKWsyQzFNVo9eT9+xIBh9cvLdf4HQVKYjc5k7fTl+cLVqVU3VoAZi+
lOA6FKODB6O7foD2pp1Va0UVvbxl+amtGm2GiWj1sfk8ylfo2hXcn/VcE/odRmRsANayZTs9zpJd
bISNy3nsRZAjPgY2/+QpsM54d3gqGWGgKisKZt21h8vjh1LULiZ0xqTQteJRqrkGPAp8aV17Xt5k
ei7QTLdjcXXD96ITnRsVAFwELM533ljPK0eEfwHLmJFd0oUrtQ4LdYtU4FxbzgmwtpsTtDwUZnEt
4A5gDBamTnMsRAWNX+LAc/yi19FenbldScy+KGdQj3QjDnSIm92PEe6YH5ezJQ0q+zi6Ikz324+D
vSpWcNU5h1OvZMU0tA8eJFPR2YcZL51KIcPxYPnEllv8xP48Uwy7/UhxWrQYdT8fXPTn+ceJ9b5G
E5GRDvbUN7G8Wlac3j8TVLgUdL9ul1gk54YoM8y3N2YgEejcPIkXwN/zaVReSOvPDV39mcxU4l3v
inIMD7uLTusJFpJj3gD6JwhCSb0FmDR4FCqHK6suD2BpOHnfHsDqQxZRGD0xGljlDSHHitm+t7CC
CqP5lqq2IginVfnByfR6t2xhOZkKbN3cBDz1fpq24dROjwlWp8mbVPduJwQrfZL8x+jm0n3DBzfW
TSq/aOHh/f11SqbzJSR/4qR1KyPvbNN+clIahjfmdMaXVDMUw/NxO3MnV8+vjAa1HJVPBT0PTym/
/V0FL530p2KPCX02kExEFJOT3wkaWoVMlXB4sHXvJI51fJLS5O1qUnZ+bZLKynFXDA2OxAgxZFRZ
cmQB3Irukgm9doUJkZaObRj/TMNXVv7tHvBry2P8w1zlyDv4DfnmwyMxVOaB42dOHPzmhn4t4w7Y
joxJtvVHovt1+W/uhLsBUsIfJIRzKdKo5HcG8OoIl7qqh1ECEWCew2T0BPBIGi3B6TfnilUdDkne
y5SQwBuGu9UsASLln9RAl62E7fFLFF90qrwDK0rYRGy7UqOCgLautS5xOZ5Mj8mHXLtZRKQODwIr
DLGtzS22zMKF1+maW3Rx6KMGCM/eN7KufJ2gITjzpJ5oyL6Yg7ZM+Iy0dGNeF73k4krlip7OajlW
QflVYUhpgTi9WeJSGm02UrIIQpS8YOJPUB8MV7rl2VkGqH7WGKMvuZn+7smicGGpWy8h3fGh+ILL
M96jw3yht6JDuy1PLp4pQMdCuVv4ymCOvO0iz/WsDtYEEAhJbemtajxPjnJO73bjD0Z1POuwLx4v
zDtVVlRrJRomRmTd0kATjyLQI2yaXiWxhT5BkcALsBz+FiXcfiZF4vHfFlbIs4tFSxZoqIvVrOs9
6XMI1rJjvV10Pn093ZkQLa1skHe4I0Gbf5oMoGRXiLQUV4n564fEqQg/cBgPOoit6IOGXBD6Fyhu
dMDyCjaxUWQFE+763hzD7GzU2IyUsoLXkdPJlULrcQrB8eESKVio33ci8ls4UauTBanNGxLaxYUe
j4FK6oGKJi4RSC9p2SI4F6tnt5QoGeUD7jFc7EvMYCmtZhU9ZnuYbS+N2v/pULmftYogtP+4KT4G
5JrLhi/NmEc4iEz3x70ln0chvwhaznwkdx6f+9Q8rSFp446kt1js5N2b1dSIIK21Q+CHq73h3Ivj
gTTcYDj4xAh6jF5m2eCItdcVT/RKa3fudlx28VuwMUlRe49QEHsits04g7Ou76Qk0BQ/NFwAlSla
Dj3vmKD5vXOlkhJ/wo5a2d84Md2YQfaHPmgXOL6VQSBw0iYjHfs+kjgYcvIWyeXrI+22KFUTwEmq
938QMtiLz9LOPBuAuwY1VKN163yWmlQH4kFaoK0uN7Fpu/4MqKnUs+pxrq8m+tn9VG0akDPPvqxC
dO2wLHDZjKsemt9FajxMvnsdvzqu83ENKZ65K2dznJt1tnhw/GHMYI46TImIygNrwb171bAgZhUu
xKcvNNzeLTeY1+la6i09ivTpGvfXUieM869Qb4xTdh/WOZ1vMGvY+JGO4kLDuBR7kuoDKm86Gvtw
4yzH/2DSc4+BzKWLIzxLKrx7bAIilg9pKhWWeFP6ZBLOT3vT9gcuCLsxdJfH4GXo5v3WeZDlY0bJ
Fd1gB8C6mAI27B8D68RM9UUxj5HVVyj+E3+nYmYi4rPYQs7OCNQXbfB0/7n0pbNUoRThXxN3ZtyG
oaGEuxHUOPWUiBm86SC0yHVOxHmSRpVlpKI6E8TM93jpvdMMWQ82uLCuyX+H5cH8058mySJdkscQ
F3HTQoTCMDibJ32zE+92FsWMARQDFaTIRt8oPvOv8PLkfDeGM1v0kGgcnpKUbhQxWn5b+yJXYRzu
SWRXd9y7v8lJ9SozT161u9NpCg2cc/RAHo6kbjZsxG6KGwzW0wNAKMiYCbSoU7Z9WgYQCM5pYJQn
eSUxo5U7JKK6bzE1TzVraTLHjbpohaQXkFv8njROefIijuOmMc7/enYNpL5BgM+GGfQ+DHWbIElQ
3WuahqswEYtDmdu2iwXnBUbShRPR+xXcPROOoG9i4V/++U/7J+04DPneoZnUGsMZEw//6CNrV0Dq
i5VQI8SB55ykHG/UTuJl4XRz/xXCD4fKP+uPZTRYkSsVo4twIeOEAFJu3UJLnL3Mdd3P5vnxNuyX
JUssfehb66h6Ffzsip9jNxwfg1In7ct9eY3Gd6pG7eEQMn1mTMUKYRF9Y4+83GL65K54tYqgUcZc
nKXtu2sgFmhUlOMAm3jgGcrbYWZMgiwYGcCa77MqGSMRPzmFSMDDtIilEP5IAy8hFDS/yn+MDMpB
YKpKJUTE2artpdM8p8ejLvXgVJ+0tN8v6Y3zLyr+NJkajk9m7wBbz0gf8IZCsl0D7vqAv/tQulKf
Wtja8GjkZ4q2eTnveIzJqJWkusQsStO9MzbMEvhykH/2sm/ko9DRhyNqEASUpxGNtyXpkrTIGy04
fkfgy2yIcYS3ypD8WAou2kfjmXicDnQlD0kFjjug2NxgNdiu9mMgNyt3OTYda17l7vkTmrEawIYv
YDpnEzdY2+299lLArLXGjEUSZN6Mo9gIZvC4KVotN01+MAeULLQvpB/RCfugLr5bwcdjeCrmyasB
tShiBF6pd8Eb3g1sS3nAeAjPitXWUkiGiP4NA2LOlXMgEozlMtlv2TRfMHh56NYqO2A9bN+65/vJ
+1/sLi0f+FD9RCbhhw/qRCFJdMgkTOHdganY959a8CszJh1DWxwNQLvx91LGqyje3QQCny3zfzBA
EYprZ1vkyVvRfg87q78yTEXseq+W8vMy9cQGx6wgyUoccMWaI9QkaQg0DjTwNIn/Ev9eL8UxaRwz
FnV9qzxpQ1JTvcy7/+xfq4DFqskaoPgIqH5v40sP4QiwWW//Z5lU0T1x7j79kjVxtE8NkWlYmrzM
TWE7W7q176pNVJ1nkpUKtBHOkvJIUnwKnooN7NNkHWQ1wlpL7Z6J//hRocgFRwQ/rEGpf65sutF3
xBC1/g55p0oCvaErZ8DOwLUZDsBLknyCsDaqj3FAgJiooxDeSUTCmC8UG9bX2t/A9VkCKK+3iIrZ
wtEa4U0EPAtc4sFqY0Xe1UVuPyq/qCTVQ9Byr7oMO3jbSn1wbenAtgJYt3OLVLlipc5E3d3ilFpp
M8pImNv46zClbuEfUCOpEURgEId11CXlcrKkH5VVlSMXmfJJITUm0lQn0U3FV5qFHz2XRsXFf3Vt
MDmreIx20rgojs2lt7dzX6dNJJAKS5vc8RHnVxGPAde3RjUydD2TdlWIDbnoifSS3ilYsk4sGfMM
JCy+MbZFppATrFkCzwhBWd4NAt19pI/8OqlSaq3DpxIY+frPhaW0ccT/9b3BIs8eCw1CXYKmNaIe
klHmEnaoft9iRt2/sYblIxcV0KrkLuELgYw2Y6pkhzP33DPHH9EyVn1T0cn6XITNi579Rnc2c6JJ
y/oM8gRhjLn8mA7fgtf3LKpgyVwUoQe7wizIKFeoMzQNTJgadnQe49be+42iBMFmyyRiVzpRGyWs
PfTDPwTt7hY+wuiKejWNBQHi1qijejZ0MsKmlQYUylJaj2T7vO9Us7ItLqXSv6+l/8r6w0XSC7F2
R4oanEtB6Qp2Meph6Xbojw9GsH/0EoMhOHbTIe8maPCbgtsMdL+xWgLxm2crZO8AzPwcUcgCvQ2f
qzODBwZec2fCGZM41rbc6O1tTta5QwHoyH7NCy627Za3Wk1cZQii3ljKzV7x7HfCRxAlVC5SuvlD
NjBSaJARh0nVdW0IwLHEEO6FU6NNBXbZY7F0zUnC0+TCGtzMaptOx6KgYj47YK7pJ5yX6pk+o1Ap
i6B38age1WVG4/4FCAO0EaCK7s44yewdf3OS+yoj72wW2ANqZCQLscPbnbBU0MSRaSrFUXJc3dBU
lKMb+7vshPLvQ35+r0CBWtc/wDYBrVuY2bt1C8bN/E/8SCqAHmhPiLRLnT5dU6HPeapUtx7ZlYXE
0D/xnTKLAWQ0KgM7Hwl4o+uOVJUBcwbrpcsq3XTl+kdJ+DKUMsvvoUOc/5v+ROYAmSPUxDxk4Tb/
lcfkbT27TwBqUTUYKyCxLwESPBWHA4SC6E9JpDlobpGYTVYpDl11U72br3yuIBlsnbIS6mxxDSmw
QO5T/5ZtL54TZrl3bwqoqYO2HXC5DW7HPyxxHQKjRZW1kUjjoKDDzUrUOmuWLaCZIplsh3CqbXFJ
UplTiJroVBZps2Zei4r94GrUAWEkmj6azUynv0sHlub3Qseg+hHMr7yfJGFKTzo9Gbfi5y4exWv+
c85o8StdwFur/KTCuykCBqj+c0ztYqimVYA43zVH4TXZklfXsFH+s3RkIqnoxnFMqCRojDWXnlj1
zW7aApz9+JMO1bCqj1ueMR7FNdU5w6SczdAnCC9FOy6x2mkg1j7jfYwV9p04/KKrsKAb6jM/ZbSf
77Nk5MPx6V06SmpyVpV3MyNDF3bYa+dVstOO8yTJcq56CqSNzk1/OhSl6cN/WkjheZOjKenA1+RY
naHBDjtrn+7NW8MDPK2F5+DY/WH1GPuJqNamHTWDoCXBFeYzVFZdCTQUdshcrBRH5S7+mXDieiyM
/6+r+4whxc1DoRZCDPfyvu1tDCgGsTSEHHeHHfnHCpMhCPqNQh8eBqO1ngVSM+XVoHrF0fQy4YL/
LnkoYgmOwDJGSR5JWnu5FFTycbJp3i4Mj+mof35zUfXoG5+psGBtmX34aIRvmvgw307ITuNtkmOU
dFGdBB2yq8C5XVHKQv+4FyAisXLolumKgkwLWLwmlLHFqUIFaJo59xDFgvRP2NnFZqIBdxTvbSUt
Tgp0B010xJ3BzcR5DwGbDriLB9e6HmUoLXlTk5oE7nSHQ850fQDBiU0XNJbcF/20hhkUoMYD3UvY
jmrEl2T9VsEOhVPFangkzdGBRDSAxkW3W4/p/pFpdhkIpiAa8HR9isKhpcQgAfIjxXYdC675lZu8
bOtUyqFSQpgywbyAUB0zT8QunQcxy+pMfkiiZ3EU6eJHvjuTJtbJGSi87JHFrb+37X8tKZrNlxhp
3tehFFmNMMM3GWx+0ZUR1pEsat56c/uqBtXmEcopxnUsUipIT2djn7TB6lacK2gS7UezYjylqOAe
5hX47xnLIQc3Hnf1FdqcSQROgxrh0pMwda4og2AnfB8z8cWz8s55CLarHwJ7VOVlo/nGOslBC2oU
dgncNU0p6nKkcs0wn964LFIdt9K/EO8uiNgzmW+ioRoyf5AG+4W2cEA1UCsqDNWLxMfeg/iHUqyO
s+2hVGwtrAOv4emE4KwdvB8Bk6FyQcE+Nz/CP6G074aDi22QO0te9qZAyzQasXmLpElzql/oQ44H
N8Ox7LnknoHIA/aZaVpZ5JZim8z6Iykr+rGn1yJRKXDoIwQ4/bzJgNNdBB1VunowEy2w9jsBZ8Xz
/PWwsFns+jvCPkYYQhBdcq6ThGZDss2dyzExBjRwF5WVoOuVcPJw7q7u1BNw1WAVGsQPi2jDX7To
YCvThYHG8ktzrUP5zvk4tdrmLClQ4t9u7H/InPGPtkiakUC+pyL32wd99g1WzwRGtyPyf9Wl4Zta
fJ6wiSqSRprBRDRVnwE6pgeuxSWE5qiwqJ4i7IBwzWxbPvsnyPJTa2iZvCwsJb/1G89LBxNQdVg2
FONl44/8o7H5HJc0NwZHMRNelyUvPcEKw8bN1Qlfqn06U/UkHUWtOcNGIoF20e4yRX78tHOYriOh
KdJig/rxEkZPdMR++mKsikJ+MORhrTGHXjzkkT/nk5miT/PHwdYe3qfH5Ri9yCpA2pZTA/v8GXUn
KoF04p+eqgMlkE6Yq8iLYJPIyuJQrpoPUzKT6TkYItQjspg02Vm9Ru3Ow+QEoQwZIz+V5nIOHFNZ
eU8Xp/FK3vV6EXn2QVyo80HzA3j4VLDEzshFeOeIzw/WYBdW0kxcV+4c5r81UrROtnYh5Yflf0LY
tmEOrQPZ0FSL5vC3kzqQvcXy/FTD6zzSz1hMQYhUbii+U1nWy4fDt2XURRw9Fd2ZYSdQIqQYwE3S
G8LglFp8qM1XRZ9eOLNlBEWXUeJQTXqwFasolcsSj8CBpX40tF4kGIwEN9au1MRqHJx4Dpk0bHHl
FWrzEsAJ2k/Gyn8km91kojS/U5hMB3uGLqF8fw1D6TVB/p83yOZ0BWOplgJOc7oD60o26fTwnuWr
i98xPhx2u4msl0N91/Gm2sWkX1yKVv21FQ3wrhJVxCLxFZQV1rWIY2Wx1B84P8AG3K943wahJCuP
R2y+qCB6tg7DgGZzf8SM6nDVD4TwaOrLIjE2PhRgWbq6vP7LFx3wX0QCk7QbrSHT9kxdogNQ7cbu
I11V6IuS6735uYOYzAWkYVS/x2IqlBv3ZkIpZ8eFRix/+1Vc/7pfKiiD/VAmeli50ye/ExTPoLt2
iwRCSScqJ/BxsTrRzZmQxOLVmXo8Faw8JJUq31ub8qB1WIH8d1svabVuBKyGvlAmKQ3eWsCTFbyA
ZGZaLpYiese2sUzxx2FLlAko3uzq0vXE47Sq3/mYLcVaAGIrFbqaRTag64sDj3x1M0HF0Z/uasdo
4DS+XiATRZVHBDgxYMzm3t7TlawV9X1EPOvxOCp1b/M5JIddCyNe9bDjAkcTiFWYZ1m+EVsoG58A
+vmK1E7Dcn7g+1vVGZa42BeJuu/X36NBzbitQdZ1369J+d5q+920/oObx3gaZB1olDwNRJ7sfiyc
pPtLysKlTkPe2iyWkYNoxIgPA7jEjfI/4JtknrFG1zARqDVMWgqaBks9hNzRWqVPZcAAQg5WShEO
TB6PYRCe3zHxBlvXBJnW7NQUrSTwne6CWItaNuW2BPOS+X+u0YuXL4h34N+SaqTmFn2V+w+IyOxl
fP2nbv2wzcg8Tm8CtB01oupqyfmLGkBw+La6PTmDYAKH9z4OtTk1B9EZ2g0xejaQcYAlmONhED5I
w6FaaT29HQnJB5ZQS1KSPUi1KUadxZZFmyy8nTO1E84ix7lAoqDZEHyZG1BwBQ8BEEhnsHWLPQfu
PGjjdmM/vEZGaB12GIaLeSahA28LnQYW2cWpqAbhK1dEW6O3hCY6N9gHAaSY5fR7glxTaUZ47feu
9K94U1jnqh59eq3SAK0G3IxET0NROREv1K6kqkJPYxij8dt885id2zs8ymSOoH4D4KuO+p46fr2i
ju/xPm6FL/5EmY5JIxva9Mv616Laf2XpZpiEOcKTD5iED/f5Ksv8iXiomeYqpqgkwp1iShg9UD0p
t8kIlD1QRgsckDblS99kNDxbqrJFXEX4/XeyZ+bVr2hLbG0AHQCPJOHZtBxZ7jVlvORCuiym1ovX
V5e74aSHaLaT08afSQXpwoMxJPVRi7Beo5ILmHc9gvOnVXdbYQJrTTAbyIogzEW5XePH64qOxTTn
Rhah+Ky0h0oiX8VKAj2av8kTOH/x3oudK/C+Lr54NG9IUBMUuo6cE4qTw0QBxGG1X21jakIFYFoZ
I5ub6yIsK2q+uTD1ed4NE61/R1lMYOODE9WloCjFY7CVtO4MQRv5AngaVl9x04+lk2m13bLHUkvz
ItdwmQJQN4kEAXLQg4rwGllvvy69j5w1GbyO7Tusbe6HYG28Hf9q6PGN/QNVWQ9cYieaILB2X8fD
pOeuQWeVfL8hqMDOUWhMkvZFDOo7Nd206iOuk1P14uWR99IHGzZ3mAX/yFRONLcfMGwuLHvPe8kb
9mFnGcZcXo7o0ffagrUnlRw6jw8jeULp/fjL4VeDLa5jYJiKjYbZWnIQqnOdCB3gVi9syI5rVliE
PVulXepcU6XPDwEo0CeZTXiY+HBoeStc3Mvpo4ZG2ofBkXj76zJ4j5E3UPj97Ssw445E3kopLnv8
aTX4EeYIwcfirH7z5Xvzwvp6ivYLSaQpLyZar/QwCskkd2K1QMl+qCXETmauBkufzUbah1wk6q0Z
X2bqWbHeUDY0a0JiPXVyVjn9SsVl6PaWtLAdcGz8QHHUwNQJwEIL/onkwg/MSlHdduOHVLUPmvBw
wCR8oGi08+M4F+NJOQwkO8INPfKPeu+skxooFDV1nk8CN6252hqrHrkOYNe3qXUG+DpFeNl1sLGT
+p3a22MESNnaWb/iHf/PQYpCaSu51JEuPzO80F4oFxsRH4OTp0vgjQvwDm9WUYEbXdPbO1F1EzM4
m1kwlNaIxOQ5lpvYw0W6zSW6t69jAmJ821fuByHUs80aiBc+1YWJwqSWoQt92B7gopSIJRs2gLvJ
LXFiI7WVfjnbB8SNwzrsbjU6SqwRwOspoHy0vN3CGGW2wSjPDuXerKgpbt6IAylwpa3wTU98Bw/u
U95GpywOMnoEO3N97MG5JB03B69ObfEXyQykvFMtESUy7B0ZlW5Ke3VGZuX3sqcAaFvswUzw/m/r
Y6jZunaXifkzjwg8ZuVVJ1FqDIDXwdnWjGB74lBajUuwAIVQFPhg4gza/5EFjs4rZp9wOmbttckS
x73nNAQrl8/wf/sx1l3sTDq1eOd2R1n3hxWmLx8rcRRyId3nZ6hfYG5PoClcRfiMvthjIREMDVtl
jsS44bhDS3YBMGaf8zGxxIeKTPm3wovDgBlHXJuhHUaXB5MtwqMu18qE+alOrlKkhiGKJtm7rvsP
/lxN+w2qXv9alIOhD6NZp4kOWmkGM8zVGsajlX49UwMcSGgmWSO5l3rVdSJZsAMxKTAXHVgZdUqb
oIKZnSwuPY8I38Z0HhVE/hRiD2BS3C2vO6EKhNTvQHdJ9aNSl6AZZmBHqBS3ifOS57dfLyJMrn2k
tqGpW4HkQ1V+RMfwEq36uyn7cGXbq8KSqjzASzU05zWmMS7yxnCPX4iY/TeAqYp6clEVJ2uB3nnh
VHBWCDxAfwghBUz41XcdkFxoulQ1OtsMrdu4NiH1VwD37r2x5+UFERaWyHS/BBXzE0lLiq1jezji
VzhGDO41o1VKWuTPPzBkmb1GnBGsXJrFIjzIYG3DB4CTuxqi+YMp0oPdUOfJv/cWNwOcHOARIrAR
FzIfrTqIlCiQl0ESyGRbWjlvSGcVmIOAXSsk/MYFPioRH7XstuBRVH9cfxTyVRSod5Q4FPP/TKv5
1uoQ8tLjf5ZyzAKFiocaumqAvZw1NTaINzyC1ZsBoVCs0h2qjg9tfHDEZN1BiTGhywE68oCaI5Id
V11RvSB2ffIqPTsRvsCVy3lMQjVAbmNtS4o6VettW5K4vKjJIbrzDpCxIhKL4evMbPjrZfjyOVpD
k/hI9/G2N7YFTr044TM+IxlvzOR0yNFM16jJQO1W3RTnSWyqYgU6hBbiyNek+N4JMGIOgxBJhuRI
nmuFabu7N5+I3lE7uRyUi/8/G3i2Mzfg5iHKOLt3mjOLXRzc+lAQLNjOJykznGNT5ixavxNkoAZq
5w2adTwHEbEhAmBU37MGUDki2skorwDyTnIVRdn18YF9T7u0RvJDHWOihOuEaXXgD0cz0YoD5hZj
P/mp7D4vn8M0vy7ZwdVx+uuWxacb/C5J2Ajc13QZw1KC8uk2G9diA/oXV6iFmEFRuUX2PWtNy2K5
oQmIU+TAJq9tUr6ppQXJY/Lhtpw2madFNUXnsCI/5C2oyWXQ0uD2mfGIjKenOmBhhwbuUEjWkjfJ
OSAte3DpeXCF6U6ER/pvbuqei854r3234chteUxAQKb++K4DbIifVGMXTYlvVmT3SL/VjAubf2tT
FljQWfRnyzYXWt03SmzUabUbeX1C24fpnSA6Pm+rjDt4dCfYHioCAOMiWBvI55vWBN/fNfPNoU1x
mzpzXEuxZ4F8bApCeG94oHYzDWIn5qXzkyGe3zhzJFH8XyaaoMLSheu72if5vLh5YM0pAdSUnGFw
PpxdTwUUppF6vmrwH9Q6+tguEitWuxtDTzUlnW9P/uSKwns1adRRkQOTKrwOu85uO8PdIlUAF1jV
x3lsrC5mkEozaIhf5yzqnqMsoOah36ZSSwHTfsb5z7mL8X3v6oA0BUc1A4qnfaWbRNVBWGQmm7VM
uKONg14DF4woX50h+8GEMbhwKjsAEFMSxZiRfIM7POqAZQ7DJkJL4RuGY106pNq6BJZ2MwmDsoZ8
j2BWluuIvv3CiwHmS5eB8yztMZYVCE5v5qLr5L3Zooc3NU6xyESNE4qg1vXJpR2jZfZSG7SdeFLw
1+qtKTzjtDD+hnHWiJQHqDfi5bIzlFkVGUj76qHcZWphjTfQbJmsmplZ+3aqC+Tqbm/PKGmwFXKk
wKDBoHBpl1Q/B7ukDR9jI2WHx0Oq8hiDfYyvS3ltQx/zb5mQ1I8ROpOtgN6NX7DaMbam4IC+WoVF
XXo/boBPkPkUsRpozTEJ3GxOtsBqnIvW2p3ZhreLu0XrA2WkDhrK2vskm35MlY/DDTk+spl/vkZ9
1AWQN3aytJ529lXIa8Ghx+gsHWzxaZ4tWx13akVGUrhR2c2WagpRKLTrhEx2Zmwqzvs9lsnL0oog
hnlDHfBu8ROQlZunOtLduZOjb1u+f0eIEs9vWewuKEbCmDaAwLj8yn6HEW+R0ckR4rH3UB/I0Ev8
f2j45T865LHA9LViC9GklBDWzDgFK5+1LQSQF/HG+lzmyEZued82j0JTYjvOTdxgnAXZHuJnvIUU
JS+SNf5BnPS/9fHpyFas7lHWWMkWhrHKJqLzarMctfcD4A//q0DqrwnnhLrRpSzvFkFIpUNsMC8h
41Rct6oC5EoON+DGJFHe/2msUWDEc2TJqSlcuXeTMmw8VvXhVy3Pc5+UgXPHF2B+D0QLqXdxoVI/
HnCh2zbdchAQiMrrAIv25iunlryLKp7VvlI1OrOHPkMsdOg1k8FAzVWlQ4/2sYLyvGw6GLpVZBdb
6TnOP70e/DL77CzLRjCAh6BfaWKS06WpLKQiQzxITNvpb4gKMRCB3J1/ArfXUdokaShn6wmv6m51
0dV6U1OW1Gafnifd98PMJFqNR6ad9ByOuYHT7OHzwBpzcI4+dVOOVOq5n8fZgKiQnTjja5tKq4Rx
S5HASPVH/B7/W6MDAirxb0Xode4T5BsSCtY4KzEU96q9ymOF7pnUivPdlt3xJVPjJgimCkvFMrp1
YWfV8ZXbWt//GJb4ayKyrtivSsasVRUUYw8iJctZcd5pHywSotJp0UODhfSBbp/gzKrR03gU0hhK
/BCgCi553X8yPmXLpW0GVl4jzHlKoCIerZ78Vjuj87s9lJhDLIVm4bylQRVLmn0OCWO7ACgBxHFv
779SmYDOZK78qVCUvaORi9+cOkwkH7SFFA9R7ruIy9bo0qNRkPWgRoByI93QejAExUaYWrZMyCPT
sbNfQjqRj/yGg3v8v/yeFndiyRqMkPqANulOOiPlMV/jV3o+uYC1AtwUrGZ0mG+fqGLKRVO/AXue
ioOceqrtMrNgOR1iXuFZogsAc8AukW1yocdwJHeZYv+cy26ojEunaLmeBVsjjyiB/0CwJs4C2coO
divRTsUoocvggerdD5Iq41GuNSCBdFil8KR5Yho/ZDbdnCo/mx4Tc1hvq5V2vK+qKMOhMn7t13fb
Jz9yX92BpxvP5m9IyYVgUFD1IWN0J/S2BsV2n0iEGnmCn1ANvz3BSJOiJol0w0ycuLa7noY8xXTO
T9krLtXUTkSYcGq2jWE0FtCCYcsuqTasw8+69Wy9atyxxBgZsRHogoSImy8a0sVwSlNeMP61wkOy
O/+dD5FBnYODjFxEwkvQi1d67paR80rLAKrLnt9KeB83mKWxCeAlV+VaJg+Cu6sJzle7EsjyRHvZ
i+5s2EnB7jyzkFwUxCOx126uNPNGmh/wGdcvrQ/XnBndpPfoG+E2RjIlVSXUTYQJ2LJvgPfQJoOe
/o79fjyi6i5hQW3eKbCHtd1JJWyp//R8Kcg65e34HYk2fIN6rObakfyHM3c32pVoojx+dGJxZz4s
67P7BecmQ4vM9POLtr5Yayc3a9FB8TNXtiIN8lR+YP6roxR2KuOfnuhf0l9g20KruWkvQHbbbI8k
5Y77dKSp5fXJoZRzAbA7vKbfwmY77gd0Z2L6IrGCCqd6Aco5v/F4Db6TeOnE6udt2S16MxZfnT3g
jt/ozbytwX8eMGsi7xm6NLaq5TB3Xnae7hUriPXMS8qPELeGg4r2PhW82rMKgQA5pW3PszxVJu6y
UpsYr38XbdVXIIAX+uADpZj0hhsAgkiOrKYuZJyOwT7pIDoX/v14f38N/RVv6Mdlk72fnkZPWiXR
ViiqCdQXjr0Ip9tvo7/mIYK5WuSWcZ9jkJtzw+O77bcXqOzZ3zSb+gOo1BC2t8xaUbTp9itsXm89
EJW1NzE90NXTNW/1LIgIbFKuWEdrhc0sd6zWGxbefWcg4vKb7++9jwACmEWU8JDK9ZGBbMfeHPaE
dR7uOOgW09BCYGFqQXvxfl+D8IBoxIZ/7Cj+32p5AkUtL80jeSdz5MLCkNznQscrdVcDhM35aaYN
mLVoJoecxP+523LOCN6dWtDRPJHCQ8ZgyF7z/NOL4IhenxpJp2MjirTWYgxoqVMdMJweIrxjQSqb
KhKVz9QyINjgplUk6LNh77yVZom6OOAHEKrA2/9Pal5kC4q9IouO2LUUrVWbxyHNOUUxYs+5ejtu
DDDU2/4Z+EBJPM77rIMj99IgKfliYPT2YdFAkMUwo7C1s23QWEdywnpFOAECMNGOp7VHs1AfR2vW
MJ7rWng7r3kzzKaFTEIOalq20X1SYJWl9OKqLUJgVAjr2p9C8N0Ug1a6tkVg2eiLpOjCpsHKGDaz
jbRbVNFS/uOtzYclrnTjZSQwt5u0a/NDvMuxBonyhSVuVyZzY3I8MugLYTpMkmvNTi2h9lHF+8fC
Bpccyb7H0mprp4GwOxxWa8Gjn1vErNWyuTFtLy9Mx1Qd0ThMCAi00QGJxEtxlrUlBZ4l19OLI9F+
YhKX6epm8XgRAJMlfAtvP0ujaqSwdTuqRALGnF5Skv31Hq06gp9eJ9Bjatkhe0dTk1b73lqomR2j
9cEKwipaVN2xgl3SerW5pSmE98SGsnRWAtvH2USt/rfrP6/bE1BcG9c8bU764yuxY7EFqtZJhl5k
GyJaB9FKX6KbcZ8t8qejGEGL7zgebt3fh0e60fRCERrkOSM9mQ3HfGBWbpRhn1N91iEJV0BBKxkw
e/IKX4pVG4YYL8H4VWQvZSVvxk5Gj4Dhld/ZJbttPLKxrWpkaw9t7AJO28I89l6RLIy/tnqsnCz1
tpmB+wrEuxv1mqSJtpi8L7vjtbg5mUMtncDRbuGbJPdJw6SnIhME8JZtIMD0rhVe11m+yPJfrS06
rpBUFHrLrSCTDd12+ebvucotzW76f9eTFagjpEMjGJcn8c9VMSw60m+Z2d8emCdyr+gTQ6AJNmrJ
Fh7RkHd8W3TNugPO6WoOU95kWCCYxk58dvG/nZzk6henA1Ddjd2PiF9ubwzjtHlHzhiitRU8lqQR
GTVWgPzOIeHhh3RRCnNj31j8S7e0dHuiQcOhyckfiapV20qflHsDq0Ww4hB6SygLu/+j6U6brF6e
pPIwvEDzbmbxUZwzRBluzx04p3GFsmy6iz04JQSlVvszQQcrVViT12NPIoJEK/R2iaOAVk/rFML9
OvnqssgNRepfNOyuZE4OnzM7iZ80ZZs62Wb+BF12EpFtZTBj34sW1A2sQlMpjFksxWfUoo9l4J5Z
X4kHasEzZ+uavfQY8ZpOMI38Lc+eNbCfLSJXgYEVBJbMMpP51H7Nr95Rl2I1mVU1DCBxuFPInB07
fBq72zur+Gg086RXjdimnHoZ+th9iCvp9pe4IvCG1jfRzdYPjb+IKYXRWKiOBWkmsK8JArSJk4Jz
nFApp2PwQLdbD5uUEXv85EnsFLyvdUBqjT+LOn+VAS8QL0AixXXROsKxNdifnFFHtoELTEy3gPGz
oqfGy91+ORQNV+fK67DmAnJq0BYWA4e22cbbJtSad7E2NuspNJM1KJ/UXygEgu41ia/PUVqlfm+R
0gBxLyJwO15Tr22hv3TjLICbRdakd+cpSCvL1k/P1mgZmNgCml/ppNJOXHVTZgq/pDl1mJsJPKCn
1GSTyH0O/SCDEJFEobdDpvAcYyJcMn3IP4+5SivX4JAWFaPJeylmaeH9X2hS3FlXqDkO4PRK0NiR
6KVRO6AUip9t/DZV4OJwW1j066KRLAJl833tXXG5y3Y0TiviJjUwdsgq7XLYmnW9ewAGh3pn3Siv
AKOomh/0+yoNVpPUYun6wDa1L74oDZDMWWdzdyhpFJ8XRoeI09PGMaK0lECvdciw8VKwgmOvYjz2
am2AowXTk5RmgCFxhXAN9nGuumrj25E1jJ+RCdHuA9YhR/hKBtvcpyE77ya9zQwpez1AcFi0B22L
J1UVfhcJ5e1dgPkBE72nSFOrMWTetk5qWuUA1L08HIAXLDLRE0l4Pua8AeqlkyJkJFjXWOUfTiKh
XZJNagGGBV3je65uMHgDq9ZyXhACAHMdIVBtyH5Q2ewvXP3Q6AUsUv0aKCKK0eNd9NC7nxzlQkx/
IEXjxjfkfIW5uCyaWKxd2ULxl0xj+6qubCIuTnQhOWMvSSeudBrY5OqtSpjaqhHFBB6dgDcuLA8X
vOZbJ9pLdHz8wH/ovn43+IlXq9MZYkPmkUoTnSz+Cey3aK5VZRyVI9tPjLU1L6WiWzBH9fsA/e34
NboOljghDudGtbAmUu5RzhNbCNLE4XwuSs9QzdaWw6v+/oofwwyLwTur+1eD05/1sUdGJ6+QCiuj
E8T5UFUZwW+kYnfBVi3eeEvHn9O+/Q5Lbjh3BQyI1QZDJjC/8HAs7/LqYOdySzDVzuJYTxM35+jJ
p4sngyDvffuXlAc/BBSIqxH0BQirRQ3JqCc3KskjuInaObQ64dmM/xX4lkW36al/CrfY88B9j3bW
vGdXSsJabn++OGkmFMHvv7ZzuKKiNxOf6YDIqqXjmGxCfP1xDSDJgMTln2vyqV6p4luMS6/4IHcH
EiB2X6PZzV42Ler2EtxA6zTzCU4Gt6XhfUfM8RCeXTyuxX8Wdy+nft1LCqLYpMAChKgpKr8GHdlC
Dl2Y0g0eyAkq7bMi3cblw9IfJ2absJ5w731wMx6mDcJ16ADawMNiTwi7BSOUQ0I9AVkfvTt5EscY
tKWdOJrVMsNQgO8yuhatsV/Nf3tsZIyYU/QxQ1REQM0lpfsr2xqxINCgzyamr8Hp1AqLi4BML0gm
TumXUfooOYwiZwp6qcGTLZWCshMxxQFlT6jEr/CrTBgxLIv8b3lTt5ivDUDag6CGd7CYgGwNe2h+
x2OQgCOskiVHLSNyXxxSIVFX/uOi5rrw6QHycg50jRf99tcfmPBKcVyRS7ixL8KAeziMzMmyVPiW
3pDbaa519p9FAiMKslDNVR0uhgy3AY3ZlZPJ40UINJPTS/CRL1Dl4hklYHdPgIBQ33uGCLdBXZWC
CuAO+/65lPEEH+/TJP2q7fZgTkgmdixndXUM3uqD8tTpPrjsLfkxyXWAKvWrCq2AXJIoORSXhTUY
Gmp2loQKUyRJpn88IyvJLsj+QD9Hn0SsZDTdz9IifHsQ8f9gyxtnV/j2cbRJCfUSP/mxCguhTmjw
i5mg/lZj5bjR+HjL8Sy63oNaK21WpzjVfCatl5TpYF7N5wndZ9BGswKwJc9OFNnob3TOlOBk/+rN
sd78vqMxvFV3pV3IEfIIdLkSX+rT/DnGSJdKsFX8CldTCNruWBUklzZtHgOeW1BsE7pKisChromY
kfUGDrdUY0wv+i4uXbxpkewcx4+t1dJcbjqFWE+QZaY+6eGe5ZYjvvhCBvibUNotEFLxtk0wuQsN
3Enyx9W4RYluUpmGVe54/dc+kg4HWDBI1sVo7BmhObF8f77EZ5cqJ46o//9nuD/n+1uhuWxLtUPr
t2ZNj/bfatqhx7DehDv5m7AdZsn8b1I83xs9j3rU6iAgIH3KHNJsYtbe0cxktjBydIK3I/RsdLns
Y5vS7yb9UuQaAmiJS5HVFcXGU4r3PbF3PA8bY+augFGawh5tTkOgT42SsJIyrJ9NxacKWmKw1t0S
6DSyOVznvhJyKy6o/TEWs/hUwML7MPSxhfg+PPYh5oJv6lA60g7kNYDuE7ODyropslPx/cp3J1zc
lqKNvRP8kGeuNZ9B+D6k6sNNsLuJBdvXD6mT7lNrkOf3+J8dKX6PnzJUGUPNVi1vzxWj3irAdG1D
c9/kIGrgcu3GDuwICiypL0vzahU1BiwdZNvtA8vXUuGRSgV5bxP6xWYt7hGpBhNGYg1wozk5EaTc
krJK+FFhysXvBCp8+EXE+5uSeazoI+Jm6ETd2/du4agK6XzOAVtWxnEAqo4jiMgDYMxuFgFGy/3f
36BTzRVO/MydAmpytbXcg07ZeH7ipIBv4YkDajBY4tJ/cmzem6jlBllUS2LUYw735ie5Tuxw5r+W
lJx3q46Z8DquLApjsYKTinLDOyU9oVWDPwjAqe9KeoEAV1s9ueYB/cc8myfLtyTWEPQQaQGJq6oT
4BasCGcp6tpgdHI1V2fMew4P3hfdIAy04fL0aY9XEm38olLR8Z6hYkyGwvqz5Z4+oZCdt3n0V3Ge
gpuxwW9Lgv9FEJ0JSpwGF/DQud1kc6oC0x6U9Ri26grrHMUMc/HiJh3oqYq0T2R3HhPKE65DL7la
dowwU+6dQ1hqx5qbtvF0qv/IhsbI/kFXVWopfGCSa8wMPztwvVrjVpwOtUiZD4OmxdGQo9MiqN4h
+6ifhtMXe+HSjIBIHy6wQrvATvHny728oSbfCmZstczR/OUjv6Hh1NxSIGU5Kc/pwMi9u+RDUip4
/DRggUIoOmHdP4hHN7Bh55Kbba6euPITONYc9WAWbDVZIKHK2QgKBAhq3ShmvDObkQQOrgwJ58nA
s8B+CSPY7ktf64APkJs3clEjkAb2Z1uwMn6mFiiufw4il/G12BvjLI1jg/40MQ9aJJvvXIkejIzg
Vn2EOsZ7i64zHutmxURbGNQ5XFt2If/eedBc3qQDgFKt8rYdIUnnKTleBkEDNKA0ER8i2RqLTuD/
jRQv5IQE7jeMm1k4LAmnIFpIf8shSUXNSgBsIH2ekOfuSmd/8iK9R05V8SdNDdS6PpHGoh+vldBB
eNAI2CkMrkeH2XilERY4V6LASx3R1rVXOv67yeJ6twuqTXevSuiPBzsxwhSww5LBJ4p3VwnmdWjS
ZvwBdvbnuDYCHFxUcIJxSmeuAcZgY+OsFi3zm+dMVO3hsYDKLEvngjUWeHExQhAEy9KsUjpdB6sb
pRSHENwKHoDT3AW0ScUO/2JlPF/x96cFG5Y78HsLqTaHQtjiPas1AzMS6VZXcXgScd62pToMNUXG
8B+BW+IStBpiJq3hqf6mg2eOMR2ry/qIhiO6+ptlz3A6gm9oqHpLoSx0ZPtChq6pkDI17pCm2hPj
P18AmBe8NolddZjigIvCARI/dn8+THEflTT24ebL/dDMa+PFjwhUvkk4957w67bG9Tk7P+aKbWJn
ACYnPzpvJdD0bBd73O+79hOV4QgqBpDaYBfjPsGo38Ug6R63CbGhGn+kZPC+T8ZJSMgkaAGkBwJ+
vXd3sS/61GGPdkZjCccthugWt5b28vsaU1x4Y61/TUkTspG97J2r6QnscC7OfsytV5SomyRCsVxN
B42RHM1jFDQeXmCDaLhTFChMSCJFy4dEf73QN6mqXEZiV33uLkmFEhFxRoFmzu7JW5yiL/JbEnpU
4yNlzstsgUZE21PRUFTZHkX63lkHFu6wtbY1StSD6L4c5WWbRDa/uD0H43FeYqQTbqMFIZ3BGcSg
oZBHviJuyooFCbWKNu0DWOKjN+bjrc5Cm2KXiF1Z6I9ZeL24ypOfxf+Qc+jPSFET4d6bUWdQTuBM
BQquZ0tv8vJrpzQ93/+nGIzmjL0oOig2VJT3xlr5rYWCCvOeG2vqXSzuPFLTwxCmxz34b5S1rq4p
6+E40FDXeCXNmc9Dr24mJHRp+fDUgTgwXRUnJ5CcCBZ6gW7RB66KYRnZzdSy9vgjog7b5kzEcyee
vCG17qmPs6rIugV0QF14xkh7Kff1D6LP1Ts6XKGbGoouK2AWD03cEeJEV4YYieIB/Tclor3L/fvP
WPSl8/sAlUxhZY1s1nUu6qKuBnuujTdh6mEKdHoME5gBgthcX4WRZRoUbyDTjTKsHn6NfC2hJlpb
fPbSWA1HTPPfa+e8w5+R0JiUoyU6xqFqJm+KU7ToqDvsbn6gARgtScGWJkKRGsqgBWnBijbSIwZ+
ic7u2oUN9XtjJZjkocUrDvX71mnYSgbSvODNrwWseFt6I8sjuTv6u/vn8jLsymE/JXLcsXhg3naS
VT7EYH6QVWTOhMMdyGI2XYNJbgP1TTsX7vvDsQTjs5qsbmD8uNJ7Qrx9+KoPQyXIQWkBzIzcH9Y8
tAHjaYkNs70UfGGW3bFm3ZcD2T9D0xP3SplRFxKue/sojgpq5nZ8oyvUiLbFxP3D4eoiAhKBvHXS
8QUDGfGOxYllnNW+vLJl1JII57XonL55We2+A3LjyQNXYaTiYQ3GIeTZ9t6HkcZl2NVuyrw43D+a
N4suryNoyuVRAb/ZjijpS1OfCbOF7OxRjrRLFmpaGSEYXhihhsC4fXYkjVhnmCIIpSX+k0pWTb3/
FflVPgHt4MxeyB24mAL89jgogOpqqFIWYz83mld3+l2qPCGVjHS9tn3egTELg6146hZSXb4OLkDw
bbSBix9NiBLS9lnK+y5wQ02jS/Ka9Q5U9a1rK4xwloFDTcEEcVdqc1czfVFVByCFs3NaToD/jJ7w
SR4X/uSmI5FRLEbYhSng90qLgAWZpj0HRTOASTlxY2A/DinT4FRMtPWuZdNXKa/CbwzzC3Jf/Vwm
rSKxCmFOke/bwEpQE9OmrnGmdlZPSlUDWO+mdsASZ2cdZESD7RtpNK8k6r7e6s7i2FhNUNNfN2G0
dqBoOmkyQL4BJ3JcnA+V1WSwfR8A/W6ir/2iL7gNSCz87T3B5bYrc2Ds5ndXcvHgVQlq4ckGnPvH
Edv1sbKmgs9HyEUvFsRqFlejTiDY7TsHRL3ohI+YJl3GKtwPFxbODeVXSKEh2AwXT5WzJIYr6Qmh
RqKPUNCFLGt5Z8SwuD48cgnIY+rUaCVnJTEy46g7A7FdYOcN05ystCic+j8CICSCVmHYHeMHbKSM
N8TzSSniUZDKh+HAKxETmlZnT2qtIdyKL5XpmmbEO7M/cKCYb5/VNEFs885t08IPGQUGR4rqgbKC
Psk6NT6u6e1WpxORShNfO88q5rvSIPPpr8CnOjJClNPvl6snYoLFBKz0qsxhIDKXiMMCN2pAQhtI
2thTx0p2h9Ph88z5d4C/uX3g1yIw43CvN6t0RO3FprDG5ExLqb13mo7e4aDBU9LYjooHTDQoKznp
EhU10n8hpCXGoX259DsZJx5xtSWLJAXObQTD7hi7zZ5l6ihxmcMuN42BdUSqOd2yY+UTk5ahSRaG
sIwFaa9pmu7iG7MsVGT3HMwe4k14scV9egDP3YUdkO/eSUjb0WqLPN2tEM0CzVzbjDwtLKj3nd3C
0MtoKC1h6uMADObKgvEEs1a0+p8VszP6yQx+NPyaJHggvYiJJiAZpWXOHTpPlzXVRUJhQ/wamf5d
MChN3cENOvTNFO4p+ToHlpeGNI+b++amopBSn39RqWWde2d95gPi9ZhZ7KsBadKs+b6rLzzCe4jc
AUP9Zbqxg935fbbpeVxpOkry2LdoHJoPoVlGGSoSrA8seZwVnGXSsze0DI30+46j1BIF8h7S+4+h
MBfetS+kTMTEBifOSRNx8OYOMqYeEy35jXOj99UVGrXey5drXcLPTt0cCTObLfgF9WBq5iLZdKzp
EidonMWkGUxj6iukabglxRELCFH9DB7RTG8GLq45jlzaC/F6s5fGSwdIxUK8s6TB4tvSrqsvMMyn
RgtJPzgHjiu6JOyJCg17GLZg6xHF6fsBV7t3auHG7TRKPC2Npru1cs8+sJJt0DIu3Zzlufvazt3W
gx3SSv+56FGg0K2nrirrThzp+fqQImTB0o80irbyYcz1wLzvRT//CO3A8Metvhuu01m7H5JmoqY9
M+cpLo5l56RsX4SVQXMOEFACRuD+PLVoJUZy6eh/Je4iigkjsHr6+OdUvj7nVyjJBHT1VCyBQT+H
sJerCLPLX9tIH/20D+Zo/RHA5BeB9Z3Oe8HD51hPTRkocjh1rb5fQ5lkKxWmcyX+PaJklvNzTSh/
g4awkJBA4bIzkxn5GzQIgXMDK/WMzVAiZmKGT+Jc2FZNiGVWB7gF6zIiGfToUXeR0cNj5fe8HGOV
MUENsEAlUG5ZklMGv9onRhlVqpYaghdQwbk/PvGK9vqM2enQQ3Y9Sql/jf2G3EWT/QKOA49d86uV
nSEwaLfOhDGBY7GE3WZD2P6XrBBT8ZTw8NNwMojE30vLdc87c72KGbe6pczYMkFvyn+KGweeeYgE
SzEwGZal5IGuL3zgFAjJJ47VCsKbB+GgbBpxpTvPtYS/dM98EaQ79XKEo5z4pvGduJKOdCVjP+y8
Dy0S2cPREgQRr/GEa61aq/ycOe7Zm/PElXFLyknqORv1+Td0xczuJtATZJ8zgA3ThXBlAQGnmr/s
77Jrxzg9lIUrkwICcJrb1UQng7zUnFiqYMz5ckjPHNWFBVvEPfI4aa+ri7d0uXOMwBMT+dmc/Ilc
B44KKXtEF7HyXr2r2YfFcOKZP1FYQdmSpKXolgp3HXUHAksJrcd4u9xX75J/MzSfQMTze8t6a7RX
51WSaEYn5DOp9Hdp3XnB/048dG24Ku1fTWYK2fKha4SWEUlvbihhWpJCvmrOEUCvj2Ve9Z4UOnMD
XqlPff7cb6uSFJqqzqDMvYK2F8x/YDc+wgi6a0e8D6q9qSJo5VGx6VsaYSoxo+JbdzIbE4H0Qn1A
tIRmEr/zQYUqP1718RLHBYxJJGcS3K2nCvFsoFyeEwsQBk4yRfWd3kvQAGgQMmMpPJBzfuLVldpB
Ka95Kiz77hYjV8qH+DGlor97kVHS8FDiJ74palj+oJ0pbQgFjVIDsC9JCwIN+DyhkdGFBQrFm4Wy
Q/8zIGYjVpQA7EjrCYcS4Ikt/ctjBll6W4sIzXylFEhRQTuT6OZGn5p5IDOz/3ieIr8J3nZoZlDv
YOnd9NdFidyhNPbO/pNpRjyNrs763SePqsu0PjdFKJc+DC059JcmO+V/DU8yVfvGZjriKzK/6FPY
tRGMDP3wjGwqvUsDhE58k98PbpSGc3JOwRbbL/hwXQvfoKZQqV0nIMhngD24+JYnSW7yot1sNDRq
j2ZHWsPWdl50sLorIBbSJ+xlJmJRPJ/7rvcXpRdJ0zupe7V2tfmp09sC+TnTXgZ5ylrS9P4rKB+h
9LTG/L3PGxVBQzQEfbU8RG3IlgGb53SPlJmmkCAA0nziDYm30fIngU6sDn5SjF30xCSIYna9ZB7x
/2lQxPAvMncnS+qwBWAamQgqIwTnTdcr858g9hNFo59ki4i9N9dHdn08pS9UBd6fSmBOkRsGBU+v
JK5odTV1BEN9q5p30JcUjiDehWkAaY2Z0SWGojODfOqDzywoLy9NM2aUw222kJ0q7Ts+3we4NfW4
jvdH3dIz0BOQR11YiX0n0W/19NbOxUIK9om6hKHwwWqpP+s1ieYGLZQlxgdcO3K9B/luNh8vcM1D
xAPNTqCb4jKSXSKrFO2gWPAbi5o3fiKokq4CUBQaHaOfNHYFECPw6MKLw6bw2oUvoiaBGoPBWXr/
ipq1rRjaB5oEkrWZdEPL/hiQGJ5ZCWwtr80N7YAExEGxgrOs8ZVoDSJJq5GGWDmQWP+MPKFerfXW
tepOdek6x2tb1ULoC00OqZo5xSYXnLGvpSVngFejCNaLbyr1H3B+5sOdckCUTnI1Mxq9VX4ZzHb1
Ey8nD6d0UV8XtsUqK0QpmVV3Pi/rdEo7HEyNa/hyqmvh8aTQLX/pEGbo7cEYXSut62gQOZ3FDyku
CHG1uPLkAj5pA0PB1gZs+rXdeK6RjbfDM+niDLFpR7umdGT8v9s0NjIM3tGTm2KmjaHAWkSQhPP4
c56DUUvPc2Te3/mn+bv4m7WVSgdakRzf7FNT4kaboiDo23pmM9tqlgUyH+wUeWXJ+ZwaF7sd74TQ
5jkUW6tPxZwUaEvFamPtt1HrrPfuxMQjQGOAV2OwXIiAD156Vc0q+fUPo6JFyIKf90kjTFfQsIpR
gu5zbXR631nPkvKCoBfgJbssc6AUgnlIxwg7xMEzJ2kkeSa8nsGMadItdR2H4yOLkxL+D46WibM8
LNWXxp0R76cagiT14z46wMw+6OcXlosFFJKBrdoS+tYlpxobSPvTgN/QDNW6l3C6l1lpXlxmWGW5
t+yJbX2Kh5CyPq/etW7ms/rRppFQ4XC8UsbZoJ8LtbV9ILbQ8WV9qsaJN0errNV1y7qiDKFhAuDS
FN3/+wL8e3Ink4iO515rssYsO3qQA7L332jNfX/Yny8vidwl0NncIWxKxhIxHdiA8d2XMcrCq0Mj
Pyom7P1EWve1ha7W4qSXjZ5ND4BDr30gQZPEmqiXmulzWZGerxyc3584P1FKvlRM95koGqM6GXNP
nF4I5dK4G+DTuqHKic5/Cm9BTUSa1o6nRYlSb7vZ4YyC2FlGBZdpRi6ud9uq8ovS9xO3Mma941+u
dlLNaBzMn6Par1RLGOKRtFTHP7nsMq4nbd6HXiOUF9k6igj9Cm5TrMIV0i/+t0XxcFd1Ul++mTNC
GRQQCpmv5MGVw+dJlzeo2vhW0NQ5yy5LYzKIEkdW+DrIgQWckxYpUr+Sz8KEn0YsWNWHpKyUlNYw
xagwcv6uKT+193nF8n52Wwew8xCHaLW8tlsxk9lJgCbTYPfTSL+ERSWR/83ChGP1pQLte12GHBWk
Mi687wIb17CkEcvQWBUvbH2zsL9azN8VcXi5IuGdzlnWzL2bd8cjmmu6Lm6zhW5mDVbp1wgd4cHy
uFVE02JX/83KI/UBaWC7xNE9TgpK/POBLUuBHslf1jf7Vi4g14HQS+4hBd0dQut21XC2L7gmfdMe
4cTDbJwOvyvIL4NpZWM08qbSKvJvQlhyPXSz/QoWKUDr4NJbUpDLSsp+LEDz7wmYpc0IzE4hMkuZ
Q7/PyTMFWzquyPd3yoqR/EGaUdQrDD3KPY9UOQ2hEp2Q89jIRUlyBNGqr4nESUfApCSbv0gQyajO
O2r/eTORWdNM0Jx+GXifiM/t8Ik0fBPL4Vg7YF3ohUJc4faVF2+Vq8GaSU9qHL5hEkQT25YAAwVz
P1Fu/FCV6Z3CSISMxCWIX2/32NqoTA4AFSLfPgePM92FC3nWMTl44ONamev89BnkuEwkCPVJ0nJW
yW7FXaQMW1wrZpry81pRgxgURbTgNtCxzDAjltShjcICndPXUt0eU2puZvO7TVA5ztDdSG/+aekk
VG48Jrze+54gsBqjkLTIUpIuSuZvy8OK/KuD093ACBP31lAkGVjr3nLmrqEUodMLUdW0T8zi/P/8
NmZq6hV2ULGi40zhaz2f8s+P14hkMG+fJXaKlDFo20kHwtzVkyuQ4VygFGwiKSnDnQciSB/3tixB
33zQA3m8hkFjlSeLIsdZlltdXRHaKzPwGG3y4badVdzGinTJKNhAZ37E2ftnO20Uby2Fpa2HfEi9
hPyfflao09LxvEEBNSjNEZgcYAtZE9OnHkE+eHrhN17iNlXRPLWZLFv5WDFqmDzKLByiKuaE7f+j
JpkbKr4DDZDJDp3kRG2ZRrghoIFCLd3Y/tRjCKipOgyQmfWqvrv3cGl8gvnp/USibwQ5OcFegL+5
FruVbYs/3NwiQSE16lmmRToQ6Imw+TJ8tPkp8Q7QcAmvBrZ0bgvKFX8jr0Mrx+AY95I8YFdZw0Kw
KV2ne+bRtLgS2tu9yd25zTGDEU/jpPakRigR3WOwBemtn2ZRoIB4eI8+q+d0RTBb/uIltGLPpBV/
RmXYixRtCRjCaixPGD+wjqlxGUKgs0SDy/SPKoyIZnXIjc2z68elBdHallEeBqNCURKxrP0wSbw9
I9mH9KC1whCI9v+u6aKYUpd2v33zcunuxSdfyHLc6PJ833XzM0iGSMbpO+W86jzu1Q5BNTvRNYwJ
dolldNaEtm8AlU4Sr7JfdIKGhZHMFtvB1Vlw/R0S8kdD/Eu4TQKPJdOFEy04wm0klD0/cBdRU5C4
iLKveF0e9dvwuzbwQ+fU/+Pso0IWv0MvzXbJIqGDPOo3wK+uMJP3m0JniSR+CeJvfqtOEzF6JsHC
LhbuooaoLnJHoTyCQkzZH2j0Qt7TUvtkC7B51aSQ9mYYNRDBdwwYU1cN1/Qo9a78c3dXXhN6ILdj
VetXzT2NjHPZQ4FQBEpf8OEcdMpolt8PYmdST4Cp1KDI/cS6N3CiIc9SJvW5C/fsUtSO2uZVW9eh
BNysmUTBZb6jNpOComzs1GMKXWZ9nOvCP/v+aJz8+OEuxTYITOaXht/5750uFSQF7xp/D9NV0MyI
iC7jm7M80AyI9KegOtFIOenbnSospmpIXyFTB98wyyXkoUtx8L2btY2q4f9UR50y0FNNytJl9ljD
HqZ3uHNJI07a8XA5sSP4HoIpmUsJupJSfu4CYBXxYo+f3H+X0SvpXvSEqkXcoW46RbvTrUnJTYH9
g9hzaYUOwMbI+c3OWYKLwlrTaYyxbQQAaJESq465AHoDGjZWOKk2eajF/dQxoCf++9nIl9kSeWM9
fI+0XQ7MZfmPxKBEYz6CorWisGUjkwjqOjVBH5DDPjcrmsU3xe6PFswDPP0scgdOMEgJoneoB/hr
gFBGotsTL/JmzfAkvr/hdOMvjGdkow+DDRnZk+AdP2rch58sMKCrwFDyA6tqM8MWQ/nffY6BmWH4
/AKSLDZmklzH1TpJLZ/SrX8Y1weQex5NqLvVoV6tHMw1i/XJ6OYcM34O6a4b+UfSRV3oE3PqogF0
MI3Eb5JDzfmg689llB1Aif+9huokqmlZJBH30OCjhs5hLdO5jhUDB5ZK71dGSTWCaiw/tqp+Clog
zSqkNQZxpBAGNjPUHfech9mRk9hiaKwi/IqszGVRpd1lxxVMibfo9CuvbXBsMQEjzkX/6GPlJLsy
lBE3HQcVKOx+bPTK3K1kIJ+YgC7dbLkA/UkDHIb69Jg4c4iZYAd1P9tfQ3oA+EN3d7oVGEx2F2ah
+Fp6mmBSKea6surFR2H7pI1zOrokxQ7Y1HTnLm8iyVM04XNci2JAkQGdWMdORPqcYvg6ZQXWF+2v
vAPS4nCwVTbPWOwEbLhrfEODn7ngczpMfSgOFgl0WeAvEl2K633EcykkYQUWQcEMD+vOw3GnLzl2
5Jjfbq3/aVcxDXry9PWt3rD0Uv3mvkOUSzraMMskMCFqfJv5r2zvZe1gyNiUxL103osdXw9teCdT
L2KC9SORDcKpHrm0Fcnn7AhcQlug3UuEti5vjzebrDLKHO4YPb2Vym84JuD3q+p/dTeqq1Nwz6QY
K79LF+ZYwFFbN7f5ghFC7SuJCmNTcrKUjYng3bdVN7So6y3FH7OUPa8DC/NWoUCglYlO1C+6iKxC
SIOSQYaCfbqD81R/7MfI0zOPT80aqFrK2yCiZB5zXv8ZqlE6wvJEl5F2abLxCAGCACP0tS/YKV3L
5tkGQfnFV8UuFxR2+da0vrbRbYJSlG+y5Z1Q8BQfE0uj7HaRlcRmNDjCTgHtApYpYqeJKY2Jp7x9
1+DJW7i6TSU5XK3G4fMwYjyXtqxEDeGwyznthQWy7JNajgw7c5uE0gLB6HrvEfWXNxQzVMCnBSFM
HRl47H9F8t/Mo/hS/m2AN1r8ogcGQhKGtpcoLMvOoIWqnL0KHmSxlZuVfJMy8E5EHf5CmOPkIm34
CM7xu91Sh3LQQL41weSBaledqMY9sS5RtHwekij/ajkpuB/6d2EV83D24YgJri+WCv6ZtVxqzBbW
L4Ro5MB6Exs1ZAG9Xi8DtElgl+nfY7jRLxjwuaWEmIuuLqnVQXQPVfx+ixN4PnrseRGzJAHrzZTr
xYYrAygtWbouxpNQ5TNnIyOqslyVzLyUoMAHotfvnpFctS2G4Mh9NkaaShKk63vTUlC38NMmheAI
PKJ+S5V6/HYIFDfNwKifxZQgHeMeq80ZpZlsV7vwRG0WKjT13X0eJdz20+HK17WzeHx95a6KTDY2
I3c/5l61fR+nJ028BED5fLRNp59bFFjaqgd0RcdHR4bcmtea4oSW5aLf5YFxEJcoaimoPlMPvKII
iw7eY1U+3EHt7kF9hjcVHD/UoIbk5J07N6DfHg/w8GIwMWZhE5R2nfNDg/8LZO3EzJ2zJxThRQSV
MOtyakqfBDl8MaX+zAV0feEbcijRvBxDSNzzmR7mOlnoS0cgvGHuR4Nd/YaO5anHl2OhrDViedd/
NU1eJCak5C7hQIvB0TLXYkRaxRCO+ae5DQtrDTjFmX9rA5Wzd1NK/i5mVB8EnjYykwrnXbZsYBgA
+6x4LQBMrD7nHauqHbdCeh1d02A00+xN/qnqqtDI70JllgAEaxS2zpd9GepLY8dmw/FGigrMblFM
6RaxEvLJSTzVTOY9TFlAFt8kyykmoDiqG4qUx3C9Coil2T//YrfOdapa3xpUv4STft8R0jf6/A83
n4zZNU/zQW3eLFPlV5/mNQLXy09gkKPII6a3Lf1n0lLceiexWLUEWPSB9pNyqv132VFTpJgH7+/T
mtJDSFB8MrsRVnjk+4ulzWWAqdOK728DB7aYNQ9lNHv7qPMfnC/QVFSimhMAhv5YjVUcTtjaCL9z
IwOXzQK9X6iIZdI21exgNMJPa9I8+bv7zzd4YfQ20skcf5fWxCz1cixQ6+C/22J81CdSlqikbGyh
/Ltsaezspym8ILmPp9fko3UFfmaW6/pqMeXOW0ejlvEjxiTKYTzfHHqGc7i2mN9wM1cNNgvGveIo
OViRXeJyT+WNoubIx0cqetwpCIuxCO55YXq+pubN19O4jca0aSZMfRKhXs9baoAEiXSJ/NkRhfdr
zoyNC0KF8LURZeYxgkEgYslZLlQI3xNMj8B8IVzqhm3Qq+7E3CGFYbJEy8bR8qE8ti+PUrr+7d5J
1qJPVgS815hV7aPMsFPJbxij3FlHCQvOKjZhhqATFYpoqFV06sO9/M8L68SPzkOXoHDBZPUMMuvM
CS2/WDkEHer2Vkuxt7FNHdWCVqAc+XtOmi7kUXcdqy7wDLVTPxv0jxWjDZAtjRPPmqfBH2a0lf0L
sOSbGYxWbV4Qnm7ryPrAMOaP2nThK4SfT/FXKyKU5Z2cIkEQpGeUtH+ZIcqx9OdiYkF9oMPKScPg
m6PdBB6EwnesacvJzAUYfP6gcIiboP3YbiWqfB8PnEGk1wxfQQzNBJ860M1OZHV0PDhnfnRThE4E
nxaJfH2UO9tPOesZv7O5vqHyoCCWGDqCvJisURgxi8fgNPtRPrI2zf6ef6zwq1kvAG0zkjm0aSAB
AK60LpcTesxr2ypQd6L88s1qxrJY6dHyZJ9NR10SBf0bxiIssQdkS3JXxWKKQQDAEFMwTSCqx2ps
PUu6N+hoUQ06ELkbU3H5W/+4IB892XxL29A7pO7OSR2jiQ0PWKUdIk0SDFm/0AIBc2vFShOd5idG
H6AntIaxcFQUxPj08c7Mc8rdQR8+9oOTxCbbzP2ZQdiqu1RBBCSatrQs78swTWuquTpvV5FNnf+Y
zPKq0iXa9gUUfla8DCvPzW6spkJla4Va3dVz5EBlrGe1wdVpcBIZRGORfnONfpi0CfsIb1wznc4z
m6O2r36jWyIkHr0l9WbQQOW4ECG6jp3SjIW0gvrweT1aGHSWPeepPTGNT5wTplDztPIsPyFFly+x
Gabv/3OZDsBzskMLfMA7XrM25DwjrxPiL/hLlmFEjgX48xap3IKjLsvdZ20/A20OnRrfuHT6EY87
Eo4SILJQY+/eZFyJ64MXeHTd+K54bAQhhuk4mg7ye4y4z+3eBodwzzfdTuvpgDpN3XUwVDhzPxtM
WDNe4qUhhKucaFoDaF5IrO4efXAlGuYQVF71nJFsVtQHh/yJBYwwlKaRK6oReNfeQR2XDsUzxITY
mwzHCjLuR8jbbHt/YZY/BFI5hxoFevxzsmiDrc1OKYOqH/ASpWpD+XYOoQbXxBIndsjr9an6xwJ5
50sXbWFrDzfEwk6jDUKpcdlH7v92+hCQVawLw9I0FAud6wz73oHchMKngJA9ApaH+BHz7ZRHikMB
gSE8dRWXRRH/8fBhSFYZBV9DgFc3zXmGBgIOa8zruxJUYo9WBcyE/NU2TyQvNpZi1rLUQ784txSF
aLAPolkaM/e4csnt668Vsf3PKpEWFuQW+HU/8je+cjyP9XIv70pBz338U4YXkUODgYkhyUVQ3G5/
JmkfqUjM7IosieRDV2PAEFQ6k1cJwQiUSENNLBB5LD5UBbDNtPV/4jibixuuk8gTdsXBs5wWL3qe
WdjFKu9uNFO7MrbbD3stl+uZW9oJDIQBqiXtuAomXLo3hnGUrQZu31W3P7hhekyUI5I+y48TM+K7
EUKHzILfCRlKEtdapL9dE5VzdrDRifHSe+Xwnt2PytLB3m4eDLZYp+Jbwl6lqy/Q4tgQRbO3P1mI
ip3wLR7BT5QZLFwGVqXdRgxBwJL1tkfhvF0uDQYCk29XCEKb0hprcTQWieuKG8+4JxoT5fv+gc6j
Mg936E+t0iy4OjTtTvWxUudS8aVWz+BxcGjcxMAB9fiEsTAoTp3Us/qnbs5tqtpZ+Eoi3E1Xjzm/
Ojq7r6o7oRLz8+EJwO2nJXl7l6zOvkDI1fXg1omb2ieRKedNnJ05CSXxoh869aegbm+6nGabEuab
TkLEw1alyUPTJs1Rtq0Els5mMYvQ2TYkQGV+eNTpP96/n8TD77HeK+hMBofQ8wittfooD1YRlbBH
LRV4757N000i4NvvVkbhTwCUXvCKozmPfVs9GWxXGrFu3EwNUhSIQtSstJbt2KQ/jfsym0rLaj3x
F7thYdFF5RzHe7mSnrdiuqtyDGDIyaDUR3VLspTylDNB95mNkmQ29B0vc8p7BYHh6VEXgb3uzJAL
0vIz3Kq5XXdArNrdqU2y8byrI2Gd757Z3C4ddsrIbzUL/zFYKrWnzxzfWu8jt16kyZe29tj/Zj5R
i+yQTO050Dz26vTCrzhSd4hXXdnSOjNxF/YPTjmlQ1q5/dJAV3RkSgHgUHLSeKbiUT9Dpa4hYNij
7/Zwn+CFx+q/ReFbTs0SmsB9mzckbCS0w6HSYehDfp6kww6axsk7p3hkaK9w81fAdEI0UWTitTTW
zloLOy09G0B+eMxrwx3JVYWSHyKkWzo1hpf1GCBm/r2/2yxq2q2Yhjc/XKpOFyiJAQ4j5L/ddkkX
JPTluR/mrHXzBG41fknWCzJhEO4YLhBkpbVtazOAdfR8jJDGgZkLRdHAEC39ZP2OAF59Bg2UO8/H
vpRGIWLua7JESBZO4VKLb2OH2FUrrY1w+Ancy96ZqbXCQ7QI42FfpMu98OPX5ZBXU6O/RSkcAUpu
JMH9BGv00SQ06USE1qNkHFsTER7CSsSPs6ehg0FjHXSe1YX6N05QszSQuqMHNOBfFH1wI9ZfaprM
MYS1/YloTnC+iNTWv3D2XYrLcZZQ4ywoOdM9anUAU0G5d4UAKt3YnazWMPzUe1V8AJz53VZhfTeL
AoG3X4BYJ6vu2DEqKKtyFDtSiOoD3KD0PcMQiWPRRFyzF+pqkLra5jUBk7amXEF6jXvkkFMlB4MN
BcrWJKYwOdJIbzl8zBbM+U2/KSB0o1/c7YuI0NPC/DMobd+HltlwPXpEPnKiE0jJMZplYZGSM1Ya
gnNM4zRF6dxMcMag80CLFNVfhCqGZIqyYmmz2aAiXvsssLQD2d8h2tvjIfcbx8sCtaJPsboQ4Ona
zsTAPlcsduubbR0zmXg/HJUQOlAbtbM9T9x5Mn3+vigCCv4OxfFmGaPikeEslJLWTsRvVjHKVjcw
S0nJ5Vq/G3yygyHlF6XQRRKnq/3Wr1lRsmeZIoUHKDHGF9S++iOSriIk+D9VCufJjkICln7bc0/N
i2HnOi2bCfmszbFTi72bYOoz3FLM/oZBP8tRDo1HVSGJdDpWVFKxuTc114CgMkK8gURTW60FEa0r
lg3ujKb6sACmqho0KSlinGOpooy97KIB/xLiTjPck9YulM4qmP/P8wNzfBXbAf6nHZ5aBC76RYwr
QPxBIhDIRdcPl+kpJ4Osu08Hkj52EolAY/545Lq8eguW2xARGbn8jwM8imv3/KwfFI/q3HA+Y031
a3BtAG4/3CClbHp1LFl2llIMHFLj/4I3k+JTp/8qCmKIaYdr0by4kHbbAKlMEHNF9SXdGl+qPCI5
/g59RGGuuZGXLAbN0V+RAKreU1dKWRwOkXHbYxo/SmjTik2r8lVRZIqgMKjVgaz9+hb/mSo9DplG
487npOBfMsv5qX/xrv4RyhIEqPSPgx/URBaoT2YaQ+Io67BiWjemiy1H8mG5FtJBMDLd5Au5OKeU
Q+6/Mmr9dzXyxH5vvLrxwGxZs/yPtJIZTAQ6XOkWTuie1pKnnn2bgEhnhkgR54yeH9eAXlVYKW7d
vGsd18yfpEv8fd+0ojRnVTJm7AVCUXvhRX89u8Kko/egmQTKlgbZMgzyaDT72MfiTx0eiYQyZzY/
jYhPrupsljZp47Q/0KbMOJoqxavs/Mu3Gl6M0zfRa/vykvgL/exE3jD2xHq4f1iJI3FE7liClg10
tQ3YQPWOAox1br2yjuh3WT8m4Y7T+e6Sr+GWtS3qEPc6pt9Cz3+TBDEV6JhmI/uaKTeF8gyQZDjG
xPqIg79op1G2xA7hVIC0RbKrN0oID4TQ/aKsGUngd3mmGxjsA0Fz2oPfWOaA5TQpjG7tvufcl8vE
JNI6Dy5CpiPQzsfkbSVy1sCcuKgIbqbm1fEPm/bLo+bXGMIzgai+WrhSScVmztuW0fha85lbyq/2
RuSYvSVPzbi1poHilRQEAkjiKeoMZFhaw+jD4aOMlv7C3ecT1DqTu2BOOQmX81l6LDbzQ9nUDxTM
S2dOW3M8tHwHRbH4IArRiE2aFE3X5G/CKfdlIETdznuhLAaDfEpyao1UNpaRvahZhzhyTtphc3WN
TWOAntXQdo3k5h7/r4SUu0gOPOai1+u+n2HH65lT1B1lHclKC2GAIPcaRv3CYz5OfRqNyFkYwezt
aS5rr/I+YoSRdcpjyLuh1o7v45KmbHzw08CRbsA9lyLUvUNsb4HxtQUW8CvhtsJoxY/uV+bkiTQa
VTY35oU6mZQicCR70kLGL9vfaVCsvoz7Ya5vUXiM9j5H9/lAIaJWiGalp9K2ZqmQWjPWXyS7llf5
MNiGJRSjf8p4iqobfNgfms5T/fdfFckHdRTOOzu2Znss4u++pFy34R+mB4DcBMhXDXnB/OBzWX3V
h75smTZZAGVzD7RdYnMfbnSGyRJ/wFv87QRfok9eQHrvIyO55FDFY3ChHXt1dsRtagVLHXPKaBtd
VlDJf1CnnLx8lxM95xapHzSibTP72VUM1ogCRdTnp4GUQVUcXxGx3lFMcLW+kNRDVqzsfaQlGliA
91XY2LiSQ96fLv7hEIkaPn1haTd3T4AEKI6KK/K5wtLaJsdPSfSjfCd0/HF2WEhr488nJUy9C97c
9LHP/HlZD1leUi890lMydL27bqzhPZ0K0gOXO7r0bgZOY/wJMcjG5a1pdtJHEwmAd3xYNsuzsvFo
WXK3zsxeRK/rfl4Vd6+zmSMz/CF02an9gMBrAVGeWrtR0xSLuj1qbESIrbeRX1lS+6vRTGMljzOh
2ArjLQlOGYb52kLYxq19NFyEykC3GoDX2ea/cGRaIWesBiXAJVYia+wKzlvDJik/zKoqdHuO11IJ
6FedliCouBRyPilnWPuku9djvFgg5a4yFtlHVVRoWcG881hxvkgBP94M9x5RbgG12cPPUGHYvz+T
w1I9OJ8Wq0/aHVGBJnhXpYTVf+LfiHj8ft/yfOtLnazDf3YRy/y60Kt7dJJs48XS2mLvlIKtbr9z
BqOjLiR2N88FDP/HiCUXUKt78qKQW9gDLkUlJPXbiHKWw6jXZxJ17QFgHPy2MMPKTaxnu/yRwIoW
nG7csOsdPg3TMNQi7IiS7IZx2w5DjgoaYKgoHomYLCYl8op/ZvK0GD7xMMBADYp3q74E+Frrgp45
ywa8tRw53pSHjjsKDiCaagcuJxmP4qjZDjKfITjJQpWhlKg2t+3pNA+m+IaBL89xN8KlRDTPdxFW
aY9hXLc6j7wdWqR400MeN6ySfQtkApKQG7awYNTyQaSvOG8QW8o3KalJtQph4I4d1PyrvgAuaihc
WVKPLA2SA6GuZSnWA0kZ8GR2yUuDL/kHO5zEfqIqqgdnK65oyW1096UWt3bbh5zQVQBKmzoo/cMb
oZlJCzvvUiIT6m7ILFwoA3Ro3+OI88U6Hl+BfX6n/SXrXRBaGCGwC3zEHt/D6SQzi4hcw+Ia63qF
9ldf3MD08SBknW2S12nTX7wTP+mSmueVEY53X7C314NQYxhKWvlH5juAThGTWnRNuEPxN9pV5JjJ
qEYIcMYlLbfIdm+xTH1Z+KTOi5Y0q1SSP+l81CBsL8hkj5pkUR6RYeT7vpWQvCQBbTBcW67h8OOx
ZT1Og3fjIwg8TauYb+w2W+ZduvTAu3/B2mb3IKx4vVm+I75Cn6yS0dmTg4dAtvIC5nQ9svZgK91W
09n1dYjih/96xxDLhK3MvUEPwmkophO3G93c8+SJbfKFn7XKm9551v5tGgeS/KDZU4nC4yfc66Lf
/E4Z2+5F5Tq6k/JZ7h4bU4KtjYptmV3i1phn6s9sB9UrTFEvX3jG8uYRTeeNpDDyeuPEh/5/xX60
AbMCB4tobTyZnLcyRcsqKbPDtIhhrSzDA7V0Wxc0VcAWcJXVXrCLj9iPbRqngeSpf+zy9jVfvxkw
8Qssd5BvzX4UpPi0SPzInO5ZOHvp4yFRYQ9ByvMyuibn/3sJCqELw5U+boJ/BEcIv1AI0rnNHrzp
+0L7b0H4bjU39DRLeWgoNsOlD3ZDVICFLitFUSNfZyaal/5HM3U3DKbFike9V3XGvqUq8IpEoLE1
J3YDH1PlkyQul2WPpA7J1SG+Ca77enNHuhxn8oh7dhbP6c12nDQocE001cXjHbAPbDUxNYhU5MPt
VdEHZKfENmcVybFH5pvNpgrazqYMQASuk+jU77bvfCaWak3rw4kKNjcUyCN5mYok8hCYY6KfLU0D
37vxE7gPy/ZuotRinAFCff8F8/0lVrfAirmoOswR31NCY3OBQ7oB6aw/H0Sn3NdNWM6nRwygyLuK
rmonE+SpjAx3+3arWhSjHCU52QbY1eshAUhBWYlLzlKgfvicXo1nPdpKIjEIVl+HhGIT+ZcWJHW5
EvxvBS9XSJ3adMmQ6mALLFkSLQzjgYm8VBu2kx/s6ymXFgK4DvvrfXmJLuTNRiQz8NBUBIq75aq2
jP1fYt4i4dvV/HqLAuPR100nBcgeqeNC8qYpgyAF4x30tZHMqEVcJ3xqf5ts5qRxYyzvtahQSKR9
0yQKV9qhqoAPufKMq+sspdNLdYPb+tNzFrWWKxyHYI2Z4Aayf9vBDGEMift7ccT95pCsMGTZx161
FytP98omrVF6/uZb0sCk+FSGpo6QkRYXcHZ8EDr85MKh2g/5e3VSlWcFV0jcbGIGQZxl7ArV4imr
FNx1yY2e1B+H62kzyMkrZ2h3ptLpFiNBpMKhWKJxcNsafwzAnhXnCMuDALqQ5Hxonh9oyPVxjEM/
qBGb0i5++FXqoVWgOvtBgKRMhfaGMZzNBjrYp2T6pdqGVWYMv30d5OO/L4vQik16vv/i9xN7fu2i
NUTZdKtzgSy48TVJVJFeNQs6o9pmpkR2C3tnwCrVzpXlLU49rT9oHGpeNKbaG/LvgOXT/aB7qmEv
bU+JycuPS7mVoGjdj7+/gqEfS7Px0xijTbnPzgCBSt22oqStL8vz4UPhBLhnyEx+I4DBX5alNcKP
zN0gCH+ReGGkRXwC0qOJfgwd1Pn9kMLPzBWW9zD8kf5rHulNEU5Kpfesk/fAyN1sjfC1UmgiV7KG
pMDwg0qcNj3Tq0uQEN0YACaF46wtQZYLW855fMR0FwCWwvES3aQna45uNPB0q/1wgp1iehiLH14t
PVwTYGmpeMvfA/LPYNU87XsiCrL7cWOzDIXODAJZhYpJGO4n3Ty2p59UKrNPrmUbBGSP+YD7MY46
zJ4NZqsSFLZgTPVPyCYN+wN7rw4lafdJ9WmIH1yI25H4wblxnX0+UgNU7DTvsxYXr4yXIVJwJLGi
Vwjklv2fg3iVLt7Yq2rzlmqqALcI/Fyg7UjXMo7hPjJI2P/I2c7DeRUOO65aBgpdCZkk1szlL9RI
DxCJHN0elbtmH/sdEChYCIrjXsu/KMxKpl6KeQ4lf6Cl2cY35/oeL5EKTBeObXAaD5+4KKQXmp7m
gOIAFAx8zAtm5sevhaxgLjIJbXbjHWA1UVlax3J9WTjOQNkgICgqEA5ljwje13bZEomK/XP02ar7
tdqZqCYkomE+Zn1OzBAuCxHSe9HOHt7aDQtgyrfN/5/+hqL8BlTBwj0ioizj1jTylFfWkupx72A1
3JcB3Qol4lngxDrPBWgurYY7Yf/RtgyrFbqD9zahIkcjMWHxMkQ/Eosz/yc4Zn/EzowVfZyrzyJk
1H8zBXCUK9O9WbTKG42Psen4u7L9z80i99Xl+Q1b5U6qJIQinZU7Q4rFvAFia6NZA1S4qOmc7bvf
yB3L/wBcAK+x7prcXNE8IHEVMJwt+Vu4cDXQhiazrYvrItoUad2HKq+x3Nhavj0//BzUjhnCcw2f
HCjgkZcHhaEmalhzOzqPFQwKk/oS+yNSF+2sE2wZ3GzGZsSTxwLCQhs3R6oeejsmA81jdfAnUgek
PrD7v002mimPiffODBVMWeiXq1aUTI2w5GhfaS9/sSLhfwyxn627yX0fOUbTMXvWl3dQgHDmG0of
plFwil/Q0Zhl5A+P+AyxgG1eXAA3gjl26dDJCoQeaFnZoR1YjHS6zqj233Jj1klWtVbtGg++dZUS
HeYs22sG62YwwLsjcse0y3Vmcgo2pzHv4Zva6e6CP/iYfDnDUMClo07P1pPm/1DnSezmcr93FcBX
vJb50kSXq6NBbh1GJaea/iHe4EovU3RPdcy7sxIeUDc/FK4dxRG2ZMH1u2Yls9lA4HXN0lGc72BT
qlEsGUpiQUBMYaleyBm3sMDZmKRyfUXxGzNSbtp7DGSxHDc7zAccyNiol5VKpI6Zi6gnwN/RBI2n
5CKD1bVtDwLe7lItEvY1KoEb1XTH28V0DNvkKZ8HjgP/6WAHpWLFdb+yolB2kpTbnT3n9IeqIWi4
3EF7g5nIHBNodKO8uKRe+3VdK2xMMVgvOuCT43QtecNeM2w0okj+3hiX9U7GuSntYf8hBXlz/CPJ
o3nz5eVomSJqtZRfvXtM3G+IlaQqzdHv/aWfBVSMe5Zsi/o/vVyfZYEx/PlLRR9sAReNgeUJdUhI
8KTwjuBLTXzHLRc7RnTZF/zIfXxunrvVzSfnAr2vPnSYRhv2gqNXD0d1yCUuxgsJgoMCfBpUENNb
pJS+IQ32NqVJGYMHBH+5dg3B9DIuGzup82XiRopy5wXyUZp0x6VReHPizRVvBVbv1P7ZxZAI0Yc1
a0T/RcA96FPq7q1qV4cJl9LTP4sI72oSozaJhMq1VfCRHPbUN4wlbEz+PSOUGlgFZcUGvXz4U86I
8T2NzJC/cSSx/2KV+SI+atkZPlPxIoFUgDb1ICutJNmf8EsKycZ14Zx739Q6akGRY5bAVxlLdDW6
4vaWCRBIPT7FlQeEkVelNSosf/pA4BRWc1LznYuL33qYXq67T1bRgnMyhDnhOu5BPa2VC2uIPEZS
j2XAHTpjqKwY8EF+dy6SE2rIEMau2LyCGmhOr8wWcdjyJEDjTWCdwXb6E1Ycvicjc9ueofSxJT7a
9aTFWaSb+IO6Ob31FQA14xpUdPke+8wopoRzJZfcnwy2O5zEfuWfyxn/CWXhJrZfumDieOK2TFrI
XEBGgeevi9pzGpZWoHhYBznFoOEGlZJYRrMcPTmPjp+RScYd9FN++MVu1jWk3OHvAstmgEjfAJoO
OJSjNoq1gIKcSu/PmNRpuYAugoem02j3Aa7x+dFG6yvRtJemSpIvNGyppT+bemYoduIbtpLlrXaO
0RSI1y0fSm/eFrZS3t2qryyN9ylhipY+WsuZczYrqgoxEHts5v9dUjwj19TtvsrgYFPWhbtBeC6N
THjhW2aSQdbic7AYTwGXy2N0BIu12bcxH8XKcgcFcN1Bm6v6pEsg03KFfoIEew9CeusV34AiY3fc
Ed94vzLcPT4XYpFdxOL1+DQTVU023YkQO2zzYIzIGVB0HLdMtKMYeP6vbWnSG+wEp/Eg5lPVEYX0
ZM06NWz9utMyQCDNrvpUX1NFZFBTRr1DyxzlwYDm453xprUDyFdwhi7UrlphcS9cH6/NvybASLVH
cgi561MarKJUb6wvssfJspZIrgpLaUNhnWmMcsHVDIzB3XezDVHhZR5PP/UBq4e/1QT8mvFRcQKS
oaRh7x/atLugjeolZ+Na+oQvBvJ2/cEmrWP+bA8MDhUEO6yRFdyIuX8rVqV3PBaCDYH5bdfm3aMD
eDPcAA/t4RuWbGIX8Uicnh4tX6UjmpWrVh+nIM0rBl9cajO18OtnKwhedE+yL6XsD0BXCkw2+OEs
J8bV99GE0o75MAbS0Z8/NLjM4TnrV78B8HmuBjThyECv7QZX4pudZ9TeP34BJSk8l9MU5ZrCVwjb
vKqiUD5xgzugowJwb4EeMNp7OomuCxcb1IyBNotvUwY3NxXV+PeqoJ8cC2YA8YeXJQhwkhlX1XI6
qY3oLaSr2yRNQOuWyxWMQcq1oeGBwllOmXrUw6WVxJ5cjoSAouYgHyZQ0C5kkd4/z5HKc1xLRnbE
UgiGOInOAnxaeqc3WnalHOGeMury675t8JeueEy5vtO2uFuiaHl5sE1Sza+w6rNFvLtwP/EsPgO3
y1d9QAfM0u7cNa6ud+5pDtdXWR8zSEbdDh8btg3ngbxQgCJ9Hczw/MLA9oFOQyS5BHoq+4TtXzNU
72Xd43fEFcUTYEUWFWhcXu9iG7YEOzfGLSbBKwYKNFt57FRidelx4E5NVGZgsrLn08o2Ukg64aud
GxdT2Dto6CFaeJl9OcQE1yv1efA1ACwfCaLOxsFKKQk+rN+2xVllzTYyiJco1d33KKpNF/oYU5Ki
KLKdkkqxd3ije/nFWoh2doe0XyEltNO30/fTac+0GPPt9J3WC1XlSaA4qbOftM3gLft7+YVYzvqh
ELnrhdGA5Epw0GAi2soxwoNyGbudEzuFGzwck27BWPkyRLk4JUhzwvQJvXqrar0lDlrFWRS2Y+v7
W32G7i3+jgDdAncU/fKB0dufn9bR+0ZTU2/amLHHEAaWDrgNKoYaJUNwhqpO9PTIFQJkKr0wMi7Z
waFR9Tkme0tehYJKThusYpkkM6hAUh9nx6tIsWIy0cpMUzOIxhd3xv+wtDKq6dkvLv/530qspmxV
W1ztPX+rPN/90sfB/e689fMdCFGEv+FIY2WVFORTxH/27HrGojViQx78xo9eSCQ7QVad0Yp8RkAS
fJZ11sqgLfyUc5aflhKwpcsMe4mDnjh3U4lq+7/wfcrSAhpn7wVEFgCj3p0j7KTo9eIw1GWY3SYV
Dr5JVvRkXHYnmr2Gu5Ky3cZp8CqOc4IfZjHOI755M/J9Xn4ex3o1UonNoBJ4G384v8j0gW8feLvr
qmVoGVFpuX++0cObqVDyYC4AriCnUpBc4psyYNtVVKOKR0RzucMvuV7wWxEIWLbyeHHLItouh6fw
1hQwiM+/WB08MXYXhXWrVo8pI9s02UFiitaSZCW7MYy1rbh/hIZNPdHgxGI1dwUBO9GTR5pbEDp3
nVS0jYIG8NuuazE1CL5sQkJspxeC+V0N48/UJ6fdJrbm86OGhaQkNkGSnqLCLYbzlzracWHvSs3w
nnmgN0NknCmcILoQjQi+R6Ts5Dh38wnC+I8HOk94PqWkYUBFHOXAX+uUSuUzEfV8AVDsFg6U5kti
8mOkrFKtjtmEvgqi6qWNqPQ47qoEmDnmaxnOTaviqLezJR7aNYA5coR6Ux4Ufj2ibXCBsIX0nUHb
77y2L49hlrPPUW5p6PFUl4yKcGnsGszqvlAscTGAVZ8qBIAYhBlhw+7X0KysvaC21ZETOCGoIybI
BSh6DzVsh3Q8NTkDT3tkbTZjiHGM1Qn8FLNFF6XcEjHB9IPw3e9jBLT4Yai2KEot8qjn4fAUmfWc
7KP39bB6DEVblyWYHNCWvxkmBvpGMmqvlRlvG90e9LCRoFEg9hJEHEtUoYQGtihCR/i+fdSIqihh
r2GYVmItMewmvBNs7anNLFfDmC6hq+WLCCWnJgynpx5mGC1DfSutIaAn3QoJHZ/oqIS6gmTb+57I
HVIKB+ZeNi+Dw9FtSK0gZ5HI5pKnJRkGvQeWCs2AiLh17JFVnriQ7uiGJ9X3cTmGf6+IkRfaP+wf
Ysggv+Nb8umHNbV4TPUgZGNkHEX1Yx3qCmSJqSBf28I0hSmvKPGJPJsNEFlKA79p1Ivk6WbsVH2Y
N640auro01O6rZJNjlqovGonaJEOysGhquDumkjLpDwAgNBgEZqoReAIUJjCGGHsMd300c5YSeqB
B6wdrAtLNkFcJ/XV9hsvmVJD1Y0BAJbfcWOquByzM13aUJfHeujTT7qfTFnlBUfhbqVLEugRITa9
+e66gemnVq0qArAkITB+F9988YFY8MZ3NOiyeV10oRZke9atQA+yQzOpF7RRhGiergoX7K8Isa+j
vOBPyFOuhfE1/2sJtObBGsPGiX7MBETfpDrKKmjaSYkSycu3LpNcNgabxij8xvyeIPxu5SFhgLoV
CAFLmyO5fYedimLF80dQ9sCqR04dD+8Awpg6aa7aCNWWucq9rmscDSdNO2iWE65xgqYh0chCv9wZ
dKDWDDDQnpMO95QRmB5TRAlcQrtktyGJW/r/9mTLZ8+861zm1ESuoAzXxQCOf0uZmQjl8RWcexF3
Cb6wSGDfDVuPkPTJSITTAks5a250NJIKiJJPnxUdf6WeUQLYJaw7syg044RRdBhljq+vSWXx3OvI
e5E3qBzhxgU3XKNTelColCrpPUE3xB44D8mTNV8OuoWlKz6EYspxkrk8WqZ3EwE5O/3mWQx4/b34
PHvI9R5HrkAAckw9fV+wQUQaHdu7R+CddcT73+8gLVHKlcvCOFdpLhKI4PDU/6Mcjz35lDGPiO26
ji2DGlG8bk1DhL7YzhwjZEmLsecgcfXvDjKrUPa1x3xU8UcGkjx9uQ4jzpzuouuDPyc8cCrgSR7+
ZKf3buQi0TafxXLIs55moTNEg5yyvWbFLTEw7ULK2/UYLtPv2g0RlreK+XBhQ+ZV6AsSec/73zHD
aTuE2lpL2MMAoWZhkUXqzCe7TjwLNMMH8e6tFMPrq73ATF2L/Lif1/k86Gj667xGYzlosrc+Y6Nn
00lQjAMvRiPOzAvgGksbD/MEFYPurm0FuESCly27z37mYTOYQoWRPgxYo3UdlQCrpm2nDgsNeRM9
Ay1M6Lv2+CgR7t8sHZfBc5aK4iXgBIqCr/yo27DjCspeBTcn4Dn1C9xZ4FCWit8+6zGmkJvnt8h3
ER3ZHiDjYOrSIhMfqbFVXZ1Nx3mEVlgH5aSI/trpwHnMLiUTxWsIbpmY6I6S2hSq9OacVX1cFi+8
pByF8ttu9+BYMrdKIIrcKbF12+P/HCWvYxrzV88G3GuJWHYudLM8A09f2ratQC3QsVSepDYe2r8F
0XeiR0fnOS92kizp1dl3f+pDHnQlOlUKiGKbpNblrw4LeHfgley7RR3jodtKdcGeenNQTT+/yAdj
qwvy6WEp+4ZgO8p5OyOf4TMdM/d3kLYDc+w5rNOjlgCk6lBVVd24URIyMDUCaYNkGgWHvxxreSO+
qjsRpPKcdDW+8IdKSqeedtygvcQL/nckuZOj6yF/t1iXIcPAdlv8LPKLbSW+VW2pv7ynp25cMxYk
eLi7cwBWP7oECLyVkZRiu6ICwXRZQhXPBVO5TV/4nahaEC/7Q7HFC0dCnHpzgohkDxqpMVwYSB/6
/BW1fWmBlsapOQfBHMjmlcJOzdAQaeuDDKy6tSunvuEAvcjezEfuZ4FGf4vzlo53gbX8yftPAGkc
6JeTykvd/QCrUt7PyCXQjAo4cnalLRPrH3XYIRjWP+XJ8PY8pdQzyDaKiTep/TYGkrcahC9BcT+u
MA3JgaPmY9A5U1acnlpV2NsGZQBZCY4e4/I0LvZdodw9VhhLGHJVHUrcJEpdm7nEgZlmaljj+GLq
X4yP71YdGl//jGDUpo9pe4FAsbLWBws7XsjwVSTIbq8WUf+COYn4iFvBuSdSjU5tOACvzgBl2NVO
8PaXWnesZoIscB1LRHI6S/tlLK9/WF8QoU7gIaarn3GQYDWduT+oaVC4fgmJBaqGFVC1EEf4aYSL
PDcXQ3cwqHiP/HfXiZsSAD6oHPCqOoyC8N50OKegks+Yr4hKrGEjgtDUzHx6vmKKtUxoeFZdsFdd
3gvtrLh8K68ruf56Ti43Bu4UGUDpjB8xvXH/UiF+2YA+TZruv9r21azi6EeReZB3SW5tsom180xW
Aiu80lxnqLkC0lSG6FY/0hqnUJfg+uWysRu2DbaKs2V0niB75aZkbCDwymrpXZqdCt80W7h2EIvh
W9xfYvyJ/+avmTPXQ+l0U/IApfx64STH25uxqonLpPrZl75XZXgWuRFhsCL2iWBP+jK238H1lI80
KWlP2BSL38oWVv1YXRGYwU+dore8qMsFRoHunKhlLJ6E7ejgxxLOubbu/2yJ+9zOeVGVfZ2Y288r
qoLTIp0ZrxhnmM2YnGs7EEGoLpB+R30eg2PahbAJLgRg8K2YdjIGTngKO+rb+Cc3HggFTiH0xD/r
35L+d5xfix5iTk5E5F1yyd2ramWfhmnPhFOhNpxbJvfX+YcQfUNe/aa4YlPkm6HK7JEVLyV7VlGM
zIoXROQSrtuJvrNVCU7pmJ2EALcAPyL5XhvsCgPlzw6vxFZRSphf5WqEu8sn5EvT1cTh/XPTbdQL
k9b6qA2LdGICCzyBlt9/MWziCCnmJbargtl+yW2IYs+FX1RQrV5Nj12N/p9NkLQP6qP7HgXU6ZfR
3qBEtYpn/6ekjBAggRDyktAt6vKb0xuBF/MXT1Dx5eUIaSi6p2Sufu9Xr+NsaVvZFZ74OFUzwWpR
/rX1AQLIZZvOzPpVn5ps7gf0bYhIl24wbO8JMzgYzc2b5nN7f+Gxi6i5nJo/2y+6Tj0Rao5qG0dg
bmqIzz+Gw2bouXP+84jrhDXCPcxjLS/zjBEOjp+vv7lL4QwbEMw1qrB2w+q9K0InOiS4mdStEUM0
38fR66g0TTST0WCb6fedJMnGNX5pIg/Vj65e/shw+L6bt4cy2gIFKRB1yABQkCdzGYXGjMDGgrdv
am+PjztWJ2kp8U60eeU5Wb9fkwzMcnRMVU0KdS/90ypnVqPkGF07AqcT3hY9rn0IvmH94qwWh0/A
k+6PUcxgL6u6126RPONS75j4OKcK5WIzAvtJdvsYPxO5cWr36VWsnPRoFquISegfAmHKSNKvlgJu
V9+5ovwOcox5EDYMUxfsQVs0plBrtXLp828qpXwVIXo245AVrcoRD4Zti7mDnWT990VXkRMndIv+
+8zihOKIOZbkypB+YG2TR6hhmLo3r0vtWMppdoVFb1kljALDTqk8PsRygrRU9S4Pb7hcdB6wxPcL
eG51O8apPGrPNccnUPD+wPtYFBw/xSOz5/fvuhl4eMZgjuabQh5uU4GobFvIKWj/aJUFL4qm2TFz
U/iktzSrElitySp2HQuweECjkVSkepM+qATF2xSnRf9fxPuNS+2TL86yGpGudV14xWVuIYQivveV
4EUQckmjl8+916Bp0V2k21H7ISy1FUY53DfJo7n4fXHwy/e28JcqU5F/ZWQ2z40oTqnNFc+FepvV
ca77Nm79rq0KU0lHflAFKNIxfKBUX7Bp70ZCSJ2hhJiFPArugIem8sU7faLYg/nOUzXZeDbtYmAp
1TuyJiFLcIygwjahKv+Y0dB1uCfRsm2z/s2mMqZbNhTwKnL0kjZDcZhUdETM9tXGtN5U5QmB2WCr
eoKpLfHJ9Nb4FB5YtQjy7y1mLSrVDJms2ceFEAdHlj5f6xxMjmKh4M0iVKLweJqTb0xp0Wp/c8HR
rWEL0JDoQk6Ckebl0sFUlizO97UCA/7JpEVY/6Sd+VdCO6AjxNHXi7VRiq26i3q6iBtXVehw4sab
AqDJLw02J1o1LQLkxnbJkoPOm75raJZbnEt8782ozaKgQ5Im0lCr1l46L6FxKECYkuwVJ00xgOr6
Ofz8vPfPfGZ4bFeeBuD2E+8sdAuLxOBhUS/fhcGkC9VBYWkqIS+PbrX2U0+35j6/zLW3RL/u1pr3
srH597XI4lDpfRGHBLoCEwbREEIHz+7/OpP1qDIRN9+Wc9r3+LD4ag9a0ZGc/kMvOAFslW0Nftta
91TQLZzsYkK5SSOOgAEtkzXBAIrNeYJ7dio4N/6h/9vjsxX2aki+wT2kji9EUm9V+KVkQSy90B7C
fvQWFiCXcuas856FPqAju10ry3qGah8HWkDgqPs7/qjZnWEYiGJ/FUGtxenhpn3kwj/GBBIeCG39
58k7+lpMangf1DvMuX+SksN7ispDo23IPK24BNcQMI1todbnuOpvxXdmqz9BNy//XTKOPMfUSz5g
969+F+bv7vraUqzA1lSuNveyXGbhJLCMRpTSLjmQ4d9b/ekBGmcjBr4UnUkbLTnPXEMe4WnUX5cU
NB1mDwJWLSaxm5HhLq/HkdP/I2KMU4LEFzJfZ7VnzEjopUQFBwhCLARC1ZsktG570EeTe+yNLRau
1b36KZATHW3fhmc7wocrGgX1nCY3N2Ng4nhmJW4K5RZD4s24bX+v2nabTTrtqqcA9cAuoEdIjkCH
5Kge40iUTh5Cx4ZGZslhFzJFc2zU0dbyCAza7Vq1t5AaEwB3vvOMMT/hJ+wevToaNZgRWcGc1GBG
Dxhm9c7607BH852ih1V2wwF8wdcsDWXWd0KcGbmAkRXz8a2OZYOk2mhaL16UsM8F11CWnek71QOq
ib9kNY2BWX84w7JOoYmnX931nLDFBn/s3b7vAlK1PMup7EjuXC1iIZqoJMslOmFlM+T08Rt6HdB6
alTxcr7HbfjpxoqQ1qTdd0Vw4jgQJHV0Q92xIKXVgrSTOuFMQZeNxeMJCPENqdToQ8Y7xUrp0tv5
WPWY6YYgGIL4TCRE8qffOg4uBsQ+FNiVePTPmsnFHPPaPES+OFkC9pVilQBoGByDPOkdgauuG05/
6aGJSnoBFvmWo6Zbc1imCCQ8pSZCtfYI1ZXNwXKbUx62/RulsPkdScTu+9hTLz6W4zpMOfCBqes9
Dq2iOTCU9SM8AFU/1J9s2bWpY1TLZR7Rosku/wpPUOTDny6s8BGinNyktQn+6Lkyhgw8fdr2SzGk
q6gEx4cBysR6UO1AESzLIryU9dBSA7iPi4FqArS8bl99DRTLYp/Zhv9RXSd7mEI9YS3ve8p8zZSF
5hQD6AT+8zKkTFjiGHwVI0U/DVUQGcQwoVk/7hHimwUwDXkVbMuI03WYU/zXHWgedTaz1TDdLhkc
tGh16ah0zWIcZqCO5A0ZTCg4Peu6ofZjzPatAvK16Tf20+w1hg0Q1fny66Te/gJLSu277CUU/jzX
0hw4tiRJltaUqv9GkgHtmJdaMmz505R+LVr9t0E6rAMMX0sBxVXLdVEG6Wx4iktot9EDZzCYokVC
ZfQTMRuL7G1gXt9wrv8szGeBjApD75dvlgtVhHvfLT8/VkqDYUw1rGgGMThpioSrY7h31LvEqjlH
uRdBk/+skYgTHKgNuq7GAqTpJDbDn3x2IujpoNnopS+st+NyipU9InckYNmyglllj8NF4SwOFAW1
3Ta3MBlEA78F0sdGZPmJN8nHnsK4ODVlfEy0l0pWPtns6aOfbFHb6wHDn85MJTmzFAjXR3h/iKY9
b+8aIa6qi5bfYkMMtcwdzFFNHgj2JW72Yi6s6gy9CPU+Bmg4O4ci2FjvFp4p5P9UfyJKR2ugK4VG
2DsvZie8AkSqa0Yl3O5g0tiHf4gyIXc3Z5WioaY7JL1pmzwg9eVzhA9Nwd1oaHvfweRrG+ip8crT
4+gEfptv4S3iRQVjMDC9xY4u/qEGIEeGy8uQ8WukjTQNPk1/7zrGgtm7Kn18sbiuzttb389C/wA2
OnUwHqyD3gz/AK8o+/juzTvi0Ba9ODSJ+ibZoFk1fj7k8qegSUopBlv0C3ZOduNdl+5w10Uhsumt
xv6DOr4kn50wzc/aavLOJMouv0HjlKOOfvgN9+W8VS5JmjCnpiaUyTK59yj7XxgdrYuuuIgW+xy1
rX0DPZPKNEQE0aOB1YjDTqW0ucnIJQVFT5dU+1IPewNwlmivTmDG0FHOcn7hOLKF2B4E9XXD2Etk
zhYDxX4xjdT+or9jpJRde7/NazWaE168X5DZHKcRmLGhi/B6QzrGXdrEpTgNC0yIihd+tBq+gR2y
tQufjs/eYaNvO/RUvDMlUn6bXZ3UaVn2/z1zTodJc9FWzh7DfT/Q6NaIz1UVo6A1yx3nQ7qyH+wb
yxIJJlakIt4edKa2/65oob6Xr2yuxr+HvyKW1L2lYFLPFSdQ5AMQokaAu0Z4ndnG/h+wLH4tWud4
gWQy77llCN7BhBG642itlrJyBcfvEvzhGn+JRAxEKJ3urAoQX3BTTJjqOd/ORQzgfIrLdd239RE4
h/rny9TFL+tcoU42nLkj8QovNX+F7LuWUE3HJAxRXkUQih3sV+krQMR1XkW7TsdQ7mGTcudNDKW5
6wzdwDw1KOgWnsPhEpHl9Ko1IYGMJojTb56NUN37VBX36XYGjxpZEM3rHQJ/HEzHghnXUi2NDxpH
U/gDLXzAwbqWAkF0zVGVLNpnANLanKsfQ18Bg0KtlHlQsltw2UHKvdEU6prAykU+0l+LNb/a2d/6
7ioheF6iS7yozAHUf64Gbf66/fQ54slWiVWG5KJlnoBCysRYEStdMjvTHqaDDTiSzHCOyjYD9qQ4
PlLJjgx/Hs9sJjxQNddGXDL+i2sRa9B3FlueE+zqGLQX4430LKx66O3nRjFbzGpm0F29uLF3O99A
UocND2QKyNiUV45AyMbrr+upCqqp/5z7R6xJAZLPvVxvP9TcBIYi7ay8OehM373IGj+llKs6blpZ
t7aSnMn/1T4ltrCM/NTZjilXVcMbXOdyedh6BBJCPDAdFjqA39r8mzNmfWwxh8Biqd/LJeNGi9pd
BZVKUTBtOHn8kUBhpf1jP/gextVve1e+7v64fh7CwZUzPahxo5012vwCtKCkDd3YjO/hroHfHyO9
XyCgxWht2A5vOe80rRSAQgiusAtlyxX/I3acr2VpwpP5jntDMf2Q2J/Lr8rQ8fYodF4G68SVrbul
QCktpsYgPxLew1WOCGf7KQUpHtZjdHO9+TBADwr1n/xl+StCzAxuy3pH2yYEHfz9+YouwyxORGUM
0tjoSqJunLoIQo2lPXz1T4GgL6kvDVFY5SG4IzJ5fyNQMYAXG8EjE0rm8EDN8Crssq017BCGLp6I
ANVCH1PnQRdQ1D5g/jSCpIi7dDEum2tocbJDKbzH7bNWxrkfH+Mt3B24cVPVRtpLF8QcJq4G5PtJ
ckdTSNIeqM3vt1I339GXgAerPM8lXJliZpYB/UXuS7Z/nMHKVUfT/MQkPrF0gcFlg3nwbKQ9HVIV
G+jfabP9YH/uPe40FKSNQCk96MwqG2SQqXSPoDxCc4MFyjz6zcuGbrsKt3uf8Os6XXCwthhGT+Tz
b3AwwmILU1nmSb9dMDBSX0rPL3UmExfUrOEivShekY+xPkb5mftgTYznnOMTKZk14O+kCHS3o1Tu
W8nUf5//kOKbo2f4VrDWagLyij2EPWKv7+NBXcZUA0elYZTydiWh14EWv7aSu6cDOth8d+VbhTvH
8mu1C2AK5RMkzX5ojkidIyM37YTW54yVIaNsRk0voKw3m4EPw3NE9IaDMyWPJlHDDyqYRnaDxqYG
bvQW8PfrmhqDhh/v5bhzdfRyOzfZZL1ObZOoyb3gK/K2fA0CkVMFWRaB7JGVqlwNB+wOPmPrZmSo
hoxKQeXfJkMWMQQ595820OLljrAm2iivZDKsEBMONJnIU5g6XG9LxtIxVWnWFF4PMaWYlVtk5YYe
oLByW9cLwMHsTP67jzu1WdUw29tFK5acjeBi5luhZPhLRxu85S8vz6/xsbZZzdC2TDqqC07Cb6cx
DeFyg7jgk1g6BUmMkcZD4WwIAYmWa6gypo1LNAxFhdL6RPEdJ64Ay2+MIpFf087tTalZTEb1+4jX
sXeDhiJ1LyWZPRCltiXLyPsT4Nf8dj0pofysp/18JW5zFHJAJwSFzvifnYneieikRkPxk/sVGcCy
smmcxU6yoMp6eIsfhwgTaGIHl5f1kVRABZnq77YkI/oMU+s2os9v4MhaRQFmRnoxkgIAJNl0buIu
wvfBVd7s9yIVhVJqdMB9W6/NEiRzPX5Plud137pRu9anMJYwSw6ZSrT405V7KoLhxXv2Z7JBoVJI
HRCs6OI61YZJ+bS1tDk4odmMJO8IVQDVcj6G8+40OsoLnZazs7I/se6ICHuM+WRPPJH5K0ZnxRYP
YUHHW0Fi1wYFC4lhPl3kiXKLRaG+wqsY7ysR2pdvGh6qt60nnk3bz9TSxOQWJtnYm1X9gyZl/mPl
Rk/IcSIQ9uMfstzJFnjYoJvT3ZHuo41oFgypX8xNkGLPI6dA+OyLmk3Po/YcgWjUaqYPkFfit+uj
V6ye2pvflOa4iKLjrY8nKDlgk034UxDk4lNJOz7XzJQR4bTvlBZfn8kxMjYoL1qbrvJkZsYxGZWB
ZmKSmy8TGlIzupISDCJLXHQEcZ0e93DR2G3LijbvSerKXXYWI1mySqyHb8MMkM0e7ooYUsfqLNOq
wUiLZy+j4/pNZPBLSlwyHPlHsKvY4a6lMU6WkTZUfyCQJ6vdSyinbUfTWVKaqyVOYBABlhcCxv74
J018sPOMHNtXCcoYqxQREVeRDIN01H151RgAmVT69ApD0EjOf67InxMYED5+5n5Al6KfS9OHo3Kq
w14a7Q4WecTP1AztO7nDXI8u9LlUtSW5jIaBMZkr7aIBeI9rqxuR/h0ksHVmWzPvmN8U8Mb/nNmO
PQtH3gmsjj24fnMedvorMa8pYK1omv8Rcr+y27Ed0Zwi8kHTLr2uFhgM53QsbqfJyFc36jtK72wh
810+KOa01JryJHeohICFs5gJpmbPci0GBSJXceeDLf2tx2aDxlz8dS5Q2DkMKn0YAAe52RHi0MIQ
ry8n0vfVEUyXEon2rV76SBN7ZvtJnyTcEuwGLAdH069Z6/1rG75awyVIyoZTgWVnM7R8rNrBbDIT
eF7Wgzn2JsK0NBAbKBAFRn9BKR2L3LRd7f0dCcU041DS+6NCSXQ6nT+MY81Rakhtxg717JuX7UGT
BOOyLJoAi+E8jRbepn8HiIX2xhf/QhiaoEqJPS39YF1Q3kqrob+qrH1pdl6Gz/L+uRP3bWOqDRlN
Ag693cgwrWtgJiT29/t57mHvtuuzN9DvZ0frtolk+3jw5wB3/s0DhmQXeUktvu1urVCqyYRWHKsu
6dRqOSfPOnKaavu6TH4h4SB+KQREgb/QvLgwIfw7VBPydo4N3IeqCg/PjlGe18k0dxXGm2X/4ccY
3MHwOGd74E1IIIU/RNGznwKB0HI0qwa2C4nZQX5x0TPj14Qs/uDMPTU9dedL6C2NcnNSBQL9rnLf
ayUxrEwoqIKvZ8isbV8+4jMe3YwqNxxQvlCbm2zuaHZtJt1jbNAEUGhl3zZi6NpKq7ekGXR0XCwU
3HSp700UvNNNanI3pxu6V3BN+c7vLaKrxJjVV5RSabm3ezzYoiTjGmFGIJ7rLSy+fHuGtIbOTBPM
ENbOlCDQyN2GvZZ03bFTqAhqaQ4jZ2w3nb7VRj9wiBYvx7idle4svyWCGqhunEY2JeU/NqdMYDvE
RTSTP5v/Vuf/pEtlPWGmuL7H5TPWGMrHUanxjVCHNxd6e/mosx0RE+b2VRrSvHUf7BiGfTjpzgPi
fpVmF2zLdcP3Mwgt5Sn+kJYb/B2T0Uyqjgm8XFzbYfKMar7+wH5DR+JPHkFQ4nxTkLcGY8LSRMHu
KJ8WJ1bn90q6b/7aGJT4kWlbFmlv8q2EcAULlliNhVKu+Xz2gZW8IkhCqW3bWfvhDqwTITFVAXde
IAs/cNMbbsrv5xOxNq8fimtKlbWikIm0DUnW3cko9jtd4BUI9gY8VqMKcqYBYrquRZ4w0BYJ4hn1
Q6bYrCi+nUZe4Xqto8wue64ehDIcDrJfc1I/wGZAvmj0jo6d/vDqktlDt5Q6+cshDMSjM2OCzRdc
UO9tuWG8qIyJdAkfEpe8XElbTf2T0L9IRDS72EJW/Mr6Vdhwkvpjd7HL3pP7YCnIuj/9Gt5ZbiQI
okGi6uevSFz40RtE2R0BjTHw7zugH5EI/dImp5cEuNK3itg5LyAA1w1YdlEEySdGn8fJ7WoPkE77
LKJ0xCNY18NIn2SSKJJ3CAQaQUQgGV4JRayuOAbOEsjMK+QMKlOFlmDtmEmfczUrSKIXkB3WUduT
hr2xWNwg5gx5AJVR1zJ3BaZlCymEGOMD7fZlpmVQRF8Q4gjhNF+Z8gxjuIhASwVQoVbg70d3I4oM
MfJs3Jd8HIiQGX3DDLb4oWPUB3s4TG0ABXvYME65BTxLns52ouoLK4kFy/cmll60ftb2U2ioQGSv
v7g0APE+bTAnM3o25VJ3WTgX1myuoJVZ2XAKLU1YeIWez6hn4ujorHWRqE6egLVtmyhcFQS8jC+O
c0L4IxLRdkfvZAKhEJS1XSn3NL6hbCrzex1b4wcpL5OAvBJAeWN1AD3rW8qCeXg5TPN+VuY0ialU
cgSe182HtkQbylb/Go69bqvYXfI5T/W3k5jPCZ0hNoGklbNGwVEfEa9o08UneyuuYhnwOGw1TWWo
eBXU7doGrEGcT/q7jh2wZN3X9CC0FN183FlzAh2uNPJiyaEDgTRwNvH5vK/V280gDpeC4NldblQn
IbFoTQxdRblptHdZkUk+HIYWiBAp98FoyhvKDQa8N5BHuMrS5zpuXb4Z7o5VEJ+48KorXdr1utV+
6615UUvOjTPaVVvHP9/ykuJ4iPPK5Ze51LdlMVQEUsMJIBBCexIwttZ1Z5Gu9pjESAriwM6fM3If
6vBw0utVeMpSL+3c/7gX1djn6wJOE8QqPmSEdFhR5V8Fqcf4SYTZ/pqbXEwFHj6vGln/AOPAMeAi
f/KXyD1UFUrf3qAlJwv0AXzU6D18Z/YFzir/2k7k/pgnEJzeHFOwJ2S0eXb3zC3ZIiMpAuO2Fgk6
JzPqcco8sTyLdkZwb9gzi8CceycgmKEkWwwXj3ZPIbtqCswvijdEjMRlRvsiqwmz07/RRlWgrFYc
jCtSwkVkhwMFCxLI4F2FMUV+l2h58tNk6MRIeKb986y41WSWwDk0dwh0FksYWXtj6+kA8dQqoVqn
1byhG9bJezgVKkwGxEUIeIDfWwsUKIAiyaywF3QO2pa4++Dz2qphDq5I96Ytr4Snlx+M9GQ0gup1
kn3mxoJIZvUtEaIsRn70jjdmtgguwgy/376qPoaT8WwDZad5ZTDz+EC8yGBAgtXl+dicGdbEDoPt
UNFc58yMv1ESCO2u5id0iB523VsYKyx1SkMJlOgIGXQ8CNvIhLup2OAEjQnMi91K/JcELfPVFhoE
ncb7PaiKRpR+9OTKW2lnHieAqjhftGY+6IOwxjBzLdHT5q5hXh7l1p0NgNb1M88KLN0AJQZmGwk9
fr+3R0Jdud6wzTSx0FHBo1cGx8M+7Va77MRfC2Lj+gICddXlTthZCJkCHVxc1Ivr0N3sNOfUBaVf
0XMD09gcGT1tIeFUVRBj6DruADb2srLqgq8YVeiG6p+1PlOMH29H4ZFATGqiO5nDux64nBRoF7T6
9ld7xmjV5NJL5J3cKPlPU8t17VALB7C1qU3hSbp95D5N8885ltygDUKwl1M1LV9/TACK2Czlmpyc
K4MULM0a6S5CKQqzntJSM1yJcllZQ4qhQTq0y6zexo4iGyEdM9Z+n9xgQdSBczzBQFl8OuX4D24/
fYIva5BNghI2WVE0sABhuLokfKru3xV02zIZ2/0alhIgW5gJ1X0r6ql+Y7ELTvF7ZsQe5rfpe5E2
RRyNaqzCoqJtLxnWTN6O6GgcZK1OSag1oMi9+E11sqIE5FBWaqQcSt466UC9dLr3pzsh9q2v6J7Q
ibkPnQdxtByWTu8cRjV906X8AftCpUjuOpm14IeR8ZJo8o12wE2BYrPlMq9V4JRABXRiEQKFmiWP
ztFcFQ0lgY5MYA9G5xHh3ZnTK97lwGrxqQhjES8gRz/xRQ+LpRXvSQ2F6scs/GdJqL1634OpQPhj
DbhO6EXnZqyfz6DLNqo5WQF70fRK8xPQzd3XDaGz+2UEOr1MVpl8nqMfg7eDIbjZ5N4auB1qEHoK
cn0SDPgE6eZolqw/Grk0yO4kumpfge2lmO4WeOJ68+6TRgDdT/FBuD1jyoOrLnhAPXjCmG+ECJLI
D0hTsbRQOrPU8QV7gIeb2Kll/ejA1dk+JX4IxHsuY+59fiPzWbpNLY9vfZR9uTRE9jCcVoOWKyYe
9Srlhixcg9QTX4ewWklebKHiey9AMmjnl9e3uxP8bYrPE8Emy2mbRQpjopC0IIQ0pL0TUAxkq/vO
l4vktEXY8F0kC7uZ6PnTLKPO1dJ3UTTh9IcG56sOsAUNLqy0oxTlfZNUV0spnJAJSeSCk91GSVDB
A81hzwgn9YA4ndXLvbHr8pHHPtAq6GhdsDae6EzyZm1CQd5RznxS7rw+lH5WHaB3LASYzYYaeS1T
X0XLQbexhtZRn/T5r9H/bzgDw8Pi29K1kO/5QVnH+ZfQ0gPhwXZxDWCQXujIHfR+0n98NdJqTWrm
GeiuVN2icRwL6cvtWVP1QujQsOoIwLqqE/v5wl9J05A0+zowlFI3Ojpyfg5mbaHssRDfkNOf6tS0
g/KsrrUbPQp6c4sIJ19sLKUFNQ7/KdURHVz3gOoSNur+/VSKYmXWWbHqbt0t5DrisqyAnraUwiZw
VuXXttba7bqOIf/c7aEmAaCMRbu+HT3QE1EdQ28ViJs3Z/0dqw4M4cd2V+UQIrL46+L3QKFztcUq
4gxm89JAj8Wb5pr4GKwGQXYi6l+jJ7fEQPL0Iif0dPQ6KkIedPboACp2syPgKLOuhBnKKIZ8KHAH
eT+PDqnYvIpV1pLZGF2d4lZHJlYXC59xDeLTgxjmH1UEnCKXb+l5hHcTK2ZLRR3ppo+keDB6KEQ9
aC9/c85Np2p4OF62uCZJlM9+TLXWXEuEsgLbROhBmYySVmPwb4t1+GjLiU6jN4oQ1K+NcVbKKjrv
5FBXzvqcpkWga3MrkpuO6fFDl96C4hVnOjm5UvduZNT563fc/G2rgnpbEVYitMisjg5umWvMlMXt
jOVk832X6xTTJ75MxVBtGUSpr07hHgRhk9YJctEl3xfD7uBYXNnesbLukUSLZeXumWQ28i/A2vvX
9FCAJJe1MasBWPtihWrE33XSzD2Du0bLOLLegQK5JKxGT+mU26bUrmirRuzsAbT+UJKFsttAYOx2
SNEST23LZOHFcCWJ1VgI3r4+MlPReNJNi++Q3tybbP4M1ucrE5mKB/Q8U8LEiZYQo+8b93gycfAd
Z8rLaHAdmGtb47pejA3ZdSpCIBnLkuW00GmMcaYQMeiTWMSKZ9QycLZi7WLIFigkR+zNcgkKtkmy
UAnU2gQCw/S8J+sMo9usqySQfe14kafC4WsoeTBbDIMYB4tUNUww5i5zJYux0e+hNuOIbPDCyO71
14QhOOgWPEM6z9LiPi0IZAA0kYUOAPAcQPzRrqaaWIVUiSwUzVIGhvICK9jJdxXmAVK1kOJhE7eX
pZZ2H3veBPWpxg4TbqM01Sbd2gYebGRWOm/qVCv6Hke9d0n7PdUhyxKOYpfKjiHfR4NQp+JPFks9
TK046zudxn+RXWG91l86Qrl4rz56+yKm44xPI+x3HU8RzGL3AEjz1GTR/fM1YETmplnq6kfI7hG5
pPzF+MYy3zM8hBH7q2J8s/NpPdqizlr/bubP4y/vmzA4BNuEtJRcJUSMljhmeVcCl8/kd9oStZ3d
1TXJSB+2PsDLJGG/n1kI08wvx57t8iJsMnICv4fFteh6N2nu0Dw8ReSRCZplEyS6M7ALqwn3lQ3p
lOHFTipYd7oDvRv3pqs5gJcJC+CDcYA11KhuEq/ixkZckoisuIMVasrKPaTijidngnJF7R//176F
hTHWP3InHwgEerGnT4hv461o6daEFoll7XYKJiiDJ6QKcBEWo2JqVXMxL1YsHBtVIoh8hZiRPxe7
MlBwfCMcC4P+URGz8fm3E6bvWT0EX94mjyKKsr+Wqt14WZ27i4EXFdEsgSls7U46fvK/Dd3tcY/c
+GsdBk9SbuAWJG4k9s1MYxr5DbMWOivMnIjlIug3xEJx6Uyi+BEQPfYv5D2Cp1TkbPGkp/P7jFjk
u6tT2XYYCkwrY9gtuJC62Fo2uvn7JnCiPXZUrU6BEu0/hbexaD9a2QjMu5oDgAMnpXPfuF0kX4b5
cEjzKh07h9Td77iAlwt2+fAC6ml36y0HSbWOcs+74waz4PwAGh5NXofHhn48sq8viERRjAjBI2FD
NWdzCyVGvngEZsv7PT0KMonbgOMP1xTfAv2Q7l2yg4WqD2NlRJnN4GQcZT7HdCLieHi/PjnkLHNE
YMWFh09csG4HzyQt//JEgC242efwgspDI7zv2yT2Pcf5r93RCAE8dgP5w6GzKtLMrIEGnynIgYbm
mbu/KzGOFQ7AhkbQ8LLA40Z2rYGLXMHsRRdCPy9FcmDq3FOTRReT1/R9c3C6Ls2tPpRAje916s0C
PdePUV6O5q6g9mUZho1kPcCzu43Yu2hbilsJBcAAob/XCPtx5C5uFSwbQGXqUhA0twRLmTwk/UXx
TSo5m58Iimjhp7JxvnTeJDQEw7V/tjfgGgGhtI1MghkNdKREcneyHFpK0WgkP54L1Hbd2Iz+7Guc
tbg+llj6/F1F0CmYWIe0IpUkxIstjXAR08+7sMAlM8Vvj48ESkrkWqDPgV27aKYBS6wLm3/TgpN/
bLXDOiIlzqg9twRwBKGnhdy13LhjM9VMpwD4rgJE6tTBwVPCQq2uLmYPoG/zNMHDMZ8CNOYsGDHj
ii9F/FUF/fvjxKFUAAktam9GwCKpcwAbJYB3K1+lTXEeac612/y3zzwWzook7rynbRHIiDW0/yhQ
Z8HwKX95LWO/pfyeTXEIsIVLHESXGlg1ut+H+YakSV/S8QmYkhG2iDg4dSFplDMp5eVt0o77+w8T
hfiy8Mok3ZdQYG63mhR7rlQieEAud/YrlxHGbmyQsPTF+H0xetILfjjhjV0f1RQ0L8j9HVQiktxw
XcUm3FbAeUqlotc0Tuh8auKCargPVkuDP9b15sEuGHXKzof4p/p7tYJXZ35D05foRCYgjBw9Wy7Z
4331oTgaROkr7iV190np6R3Bto2XFTpq7RPepigty8oXe0iK80EUPT6evndL/6fvhKQEFEl7JzJ+
m/N8Dar7TIq2uXwb5nLaJKN+TO05x6Nq3OmFpxWKXH3EjKQPwbPE+6nDxz70LUABdOP+OJRVauzV
m63E/dnGx85ILlsA0bgZnBfViV28MgMwyoY7no3RBtlCcLBI9tOJ72KkeFAOxEuz90TxZiVDQEnK
0rYnVYRUKe6OFOu6oxQVDIg61DdD9QWpFm0GJo89PuEBsZUkZ07djLzLDJXZu8dgqgI6oz0C1dQO
sVMkA5QH9L2xYyxUpP6Vm/gkXSOxJ7WtvtNaIobFIvg913rYeaupscjCsWU5MXjzLtcbE8jZC/ZH
UGkBBeGcz/B7e8VYPPBZybqFC8f+01lBLBVqr/OWu37HCBgbgXcAQrPm6R88jL0RrbEV1efulat+
FEcgIHKxpcmEDfG54AGtszys+Y0qygrpxDrlKpUOaFV98kjsF03H9eA3sIZJBpEdiu9SbPqzu2t6
D5hQ4UtKrvnvb6YsL8Agso5fNDPdqDQgTywQ+amNznylYfSjcyzlAuYvZBMr13rzHUFxQ3Jogd2w
Joa1qgjSYQMO4QZVhCCcMloFUNcpaLayZHSkJWoSIcfy3ugZ7zTeDYzAfUy60gXUMX/OamL9wXsP
DDR6yBMml8lCH8zNhFVM9SICaorVU1EP9I11wpqOeTPScVWrBJ+SLvgSlq9LOjPAXKkaBFac9ZLu
qLZQv09BvY9ZeFRJxbPrw6NRdFaNT6FN81xLHhsJ6uzbBVVXG1WVwhF2t87NjNbQWzg0l1LM/xc7
RbCyNEayeySqZd179nPRaq8Bve3u3zL3OWLDPZE6zfZ4UhzfPbxY0yINs17bCBvmiCcDupEnLoin
a/1H08iBt9DO8S5tqZMJf+930vcF3Q9WJQncOeHP3pMTezAuxxEtspiKjL2dg/vaGFaSZEQ1wvq+
UW/y2KP1V/CO/I1A/yDdSYn8p5PIpUK/6QnkTnlYQD2qMB9cVwZLim2BqrTtE65lf1Kp2FZpsW0Q
QVUliKKg1MSoxgycCgVvRw7amesVAOh1OZ2kll2MmkP/Vrsz4VGWqeJoIIhkKEkNXw06Td7ZS/GK
WL2vT69/7rq8igqQDQ6RaPxImYW5b5K/Cjya0sBJspGhoJQnQ2UNF2yTpmShoccRjEsNr0Houyu9
mm+0GzcLp4HxankP53svK/Z5YQgNPP3xG2Q2JGzcdghHOzEQlKf1Qya658NJmPil/IjSXiuaYTkp
W1ZJzGPLcMRhBD16eY/+btTaHZ5wCXZ+YoY3CSRhk2kX/ssNpE3YeN/V84KbnTG4PbW75vrGj767
UFEBXe1qwJDiJEoTBmmubKBlVQzF8ZzMiFnOeqUwsJC1eoy45O0vvvcVz/PQkLuGuckj9ciUsRcL
VYHTuTZe0GFS9UFvkeA10ROPRwUlY4vviWCb8ZtvCs3V1oKxRSW07HerXdSSWq6p/nXQRFQlWb5C
HpQmxt1+vf+12mAoM2xtQrMlvlh6qp1XEzTn8w+Pj+/gxZ9iU7YIuMim12Rk1VlRzYIN8igM6Yrf
42q1AHqw7zzbBKMj++02Sm9++UX6FLcFn6C6DSRsnfJXRi7SF6Azo4C/jbfNIr+ja21bJYhjAtd2
6aCjM+DtVN706smzCwdpqfBNpuD6N/C4ojakAs09Pc4kk6D8XY/7VU53obXNAn6eAZlmsIdlKxCS
j04NVIZE/46+uI09+J8ov+Vj4ZyeImflzF1ROl96daJYVH+sinBRtbv4h10I6LMym8hem34WR3OF
O7YfN77Xqh1whJWnSGj+1utTLsZUST+gsQ3hJ5o8D64h22MQc7PBlxwQTRN8jfrQohUmjllpEq2Q
kO4OWYv6QPVM7lKOFLJoJp8e3RRZVbSAv5f9mbfoJurNbTFqg1FP46vRRvFl/JHDvkxM38Pr1HU5
95eoiaVLCA8jVMr69KDYexl7Mv0wGbW1JqIQ4ixCOz8janYfWcdjIr94Snab22659Ys8oWzvoSO2
CsITlSIY0qZ9YEovEHvJ/IxraIx45CyM4/RN2wqJE4Pyb48WP6NhayJHJIjOdGVhUQG7zdjWWwma
ChH+zUep4mfHGBrdDsp/MkCJQpqY4rmhWGq18sAz1jtomeT1NhDF3AoJER0eQhfsDOUOQ7ICgBbW
ILr9kPos2Cf0R5s9eqABHuzq/pHciJozGQrufdZ4i0qwV9HkkeIzaUewwOE0FohGQT4MPiUZlRFw
gX0wEU5Ku9QJA6dYm4xSogEZ4qrR79sIDJQUGHo/pLO4vLMHbhikJIwb6vi6zF3nKMZWp88f05fI
zAoJ9r/IJ8qPkCeAvrC7xJqBXeb+oBibactRQ2V4sr1bpjJ7Ig73SmRiHiM94g7ESedlrhyjI9nt
4sqs4fBYiphvyVOTAG5PBbfWb33U4B8SRdkHTZfk7H1Vu7cANlTIkFbg8k/KCFriCqsrAjqVU7sC
DoJqOFn6+5NMMq3f/Pn1rFOzaiTz0zhIbEhJd0uI7o22b70v7dVpV7ZV+vXrLNFKb8L/ZzFnSXWN
rAGXPiKUeJlhZTnobSWQuLDtULW1xqFbwY/aMHFmubT+qES+SbLUCaH7d4y81I5Wibv/n7lij5L0
k627Oouramc25G6tdOHIxFvnVHvMBcQqm848dRlz5S8KPGnVRguwX4fVYeUfGhW4F6cavI2sN/B+
gJz/RSqFNc7NclJsIvzx0yU21wIXi5AHGFqUAgcgF1logZq0s3Lg11IlW+6n50QjvrpU9JhlxVWJ
oJPVtJABeE8zCeVZlnXzA/zjs0GZN1DsQjt77mB38G7H/s3aRfc/XyUf8wM8km8GhjRSVtLHSRMN
vtFuXqkS7Pu0tFjVbW7Yu5MLXlx+qDDnjHvEJKC1hrZWmUE6OX4J/YiK9BRyJYCngpl37mKyTXRp
IijBKe9qUZKLBsDjyqPg1b2Qlh585i5dTUBHBZ7uSIp86IvTe8qC4TnpQlx6UKjaC5pVEfmR3qBX
FbvU496OR91JnP/kg8AdDG5c7c8YRTPKE44/1wrklyYlZ5uTU84aY0WlHBAhvjOunUQ4K5afPssQ
7mXSjHl9JFOXPCpwEV9jA69//Je41spd93YEBMO548/FeKS3rBgiqCHsAz4+9rM2+3l54dVLOm4x
o4fv/hPZOJ8WfzjomiU0i92u58Crste/sWrku2ywKuCaTW7TF0eaWUKoUuz2QEDWWDhclOww3tvi
o9U5AwMpN5vPTbgttdtJaumIQXArLhQPzzBc7+1bxo68aA3htvz91qMsq0klc1wIWkKxEx+kexPB
XzFKZ/ngbgAowdYpeSJ753k3Cxnn4VP2k4Q8Hl942vL414p1rMLKYX8q3cerxfoS+Ybow9qchkW6
xXjnjAwDFMmHwFT3Jt3UEAPtQQVsEFw9gZ+y4uItft1vilkKf5woi4GcBfdgTkkL114u7wN+kYp2
5Mk8aSfJ4eM46aDjfdPZpCa+WgBk9HM0yiubZ5cbToHw8Z5J+G9BT3bHQyEHk3OLYrYf1+rK3F/Q
gF3JH7rR1HYt5Am2BB40YNX1rbn3RNQg5l7IKUzkhPQBtgcVNbFcl1zaFHCioGvkjmVXuS/wGENe
Ju5hXixGoMmo8Pu5FfNMKzPZ0WCrl/sskU1WhnFc7FIyyjM/BxGtVbdlRX71RyIbLBp1YEQQ53ZY
bdQ6+8M7xPD8pM7/6rvqQRd+Ow3hujU1UeXaWutirjywQ97pa5tAkNco1zxzz77wpTa1+F3uTGDA
k3LUHDPqa8sl4iPMxDbd6R7Zr8H8TAxV586Jrl+OUphnJukQs2rIYZtH94elitouQoIpLlf+xWPR
X7ONhHuCtRQhhGXO8D/fOONEN6z4yoG44e/avGw2r4KYI7v8iGXQHn5rYlJ0nowOoAWs3WwlFQoG
HiSAfyOiOwgdyxSI6cOcsJqFS8a5+9Wb2YZ5XG/+FYLWQd0am//WPtGGuX+OYB2hpe/PMOsarkFI
uSRReQwCQvQfagZdUMEQnWqT5I8pvEwGQfFZljIVcRBw8ZbqHO14Rwg3JKVtcTuBGO5oA4N9sKvx
5kYNML2TZMHe2K1ljgMocGNQkBucbI8aJVSirsMGYqV18KAnrwMVZJ9li0nshzJ8+bfhj9qrCIxn
Lum3I55tjdU3BPQekn2aQ0/w0CpLZW+6ACnZnv/xU0SVw6a4fLXP9k2Rh2JR5SkJtewOOYZ7XLiI
iv8vt5YuAtGxu7Qj0nkCWMTUPAlzIUgFB3lQmMURCx7wY1dp00gj1X+Ivr8LfMILpkqwnVBmgBGe
/gKBQAkoK9evFEJy/RXouRO0MeaJhcj4yECKLOdGXPOem93h3uRLd3HBk761Mmu3O/dTM/8qwcI+
qcjC5578kZPHB9U0jb8O4IsbqMtvQVc2UWHF2vXqAkgxnsqOu9MhAz0GngvIawIB5KCDIGs9rl9s
PnGCccH/x6mltn+l33gbfNshGL3gAtJjS4H9sg1+l8PBaC+e3JRZ9prbGjGFeUjElmE5wovtJJMu
pd2GlgYnZ5Y8qC1BQSDk7uRdRkk2MEVKYuA1lCpvRF5L+PaX1nGO1bs1spGPPWcUzoXuqIMewlif
4Al3axmxJRhQOVSM8WJ9ggrXvaXpdCcyqHqgMoOwy0DBt2YzvL4LUpHq0/c8FmEDaByT+vj5+Eqb
mTJ26xN6xGhnNlEC6UXQVNZRlbDwTmZuNyM7Y1ZrrHGhKTajbNcascSvvfxe4xPHNxW1rvuTqv4o
+LsOWeAUMFHrooG2f2ER4EUcHUR93YNoMYcNrU8CCO5+Qv+Kt5lwETES6xMmMJnyzalcyIxuSp1k
dzQIeOVJb6M2xVwn2ytjMqkpT/QIxe28uoBAQYw5h6/oihd1KBcSrFJf3XF+zQhqFlVNUZVQraaZ
lkpDdvMuCoMEsOvoRfiNEcXbnaPYs4BJ1wLwsZPKKVQVFqiMPxfloRyYkgTb7Q74+g9A+oULpJZq
cDbd0nCQvAIW3i8EVtw3DzW415H/Q6fXYDkFLjjf0kOTtMs6HjW2ZAHu9QkmDoU7qfY/ay7uHpVo
O7scamKRTC2wUBTwBK4XpinY67kyqPGPh2MbdzD0H6dRRHSaO3xuAnO/O1aDAHOc+AI4tdmJM+lK
Umq1/9BCp2SnfLJeG4Em6feSEEep69IbKiJ9zbFzP/Oky0pZq2AbWWuM+0SFz/0Ra72lvq5kaSEZ
wRpSle4Exv7+q3xHulHK7YgGumoX1NUAeFXkZqQC0pUWpXr6lORNr71ZCiGk3JxWgoVjK821NjNO
oGfRk4eM6YHVzUa69DBTiIimruHSOCFuUE4DKTw+BkxUDkVhTJitJmnSIkR9A6bzNbOy7bWP4UDy
Uu/TeRXn4o/dKQJg2IiruYbtlkgOsfUX2XFrNQmrIkojx+PAiVMsqhQOAbiBoOuGfb7fYux7UWkR
IFFGmYFGSLqUJ5ROj/V36o5Z+owjXzrlyBoyLlSvpAePNPNtRYch128l60zyckMLLz0NPPt5weS2
NpTwHHeFsOCHdPP5AJ5UBm+yieSDPwFz5HtwMjkjtX/07LTYCzlFpvJV2ftUIJslH+q+CVm5jMYU
42QY0Z/wjJ0I61uGReAvd3ZJT94C93nTeSqpoK0BAYdryuaMfdKvX3s/tCG1ep38EAWutYyWQG0J
YQtWMYbS89iDi722BE/ipUCAatzoi65ipi2uXCKoEcfxnDDZpzzQlDX6BdET0LHNNkfYdWtaq1hM
UqtJbRPFJizTEmA2s1BcXDWeZDSpir204J2I87auHTAMLgqv7yWLm/ilhuu9odtDZN8Uo4cGFBNy
/lIZ630LjiPtb0LO3b2MiRP1epJl2aE6qOrAgOQOl8+TNmGNa5XA9w6LkNbx5CG3cyHqjJ+P5pAe
Ltki/E2fPIsFNxFwxjlr9iUvUaqg3Be/VGmMMuU/HuQ2gPffbMP4HfQvVPpKmE7GW/bprzl4+gsd
mRYxojqHxsofS7MCHcmGh5Rm9x1WPs8DBKBOrq96sshYw/YLUJe3JCRVGF2cOfqnwc1htKE7VuZ9
JbJ5/1bACVwQKk77M4+JHACUbZF7JWw7fddAzUbKeWWjgMd4F824lrLnX3f/M8p0KjA7jmmJhYEc
pyZzJKFUCNqV3bMjNl7EsbE+n8EEYx45+ZnsXXGMRQgwVlxrAL0gFeZsbiOMCcBkSastAIWEc/ey
YZsdBY5RBpND0iMc8RtltvK8uNnewn84qZRYFtm6bBfiXlNHoSztEIJh9K+ggG6FOAwfoQxgvbcK
L46G8a8HTAtkZq2Uq4J2Kms9LLlSV7FS25+/q/1DU+FxLxWlFymr9q2ibD3ngK4Exsdc0hc3mbhF
Epm69BECSfk74FrekNB17PDaFiwXrc6mxHucfH1Q2SJoKDGi4vw/k4NmmKwsCEQoRNCr6Vzu34rj
OAR47+HBeWKPU00DRR4NzlGE0Z5ugASycb8EKkBBoaeRanvPpOE1PN4RfV8cZsABjW1gbrpt1d1k
WGS1IXMjhVzYZqfqFeBrngVsAsjt8f/fCWBV5hnMuWkPMKJ9sO9R0k/5XMjq33sMjKOCf3mzdmGk
xqlrWn3O45hq4UiGsZj7U+Gt1ALTPagJK2sIPv12HRXzo1UpX5B24jJ1qJoKEsQlLoqQ2J4aevtS
gEy3cSVtgrcjiJanY8BkEZoST7V9OJDo6QmlvazwSmsnZAwZ4pLqCfOsxZKJXyK91yv2V+tMve8l
IkgldqImn29KPKTrhesEVdPs3HSsFCgzsbTQkxecceh/DheeKN2241lZUGMWWCdcK2jTCDBgT3bu
H+HVvmQqfy+M+csx6zu1EstXR7Hu58ChCCz56UFkaFY2KNyprcxgAt7cSKFM6cHicnlmQ8MjupZK
bE251OLkZZiaK7D3VjORaktgz/LQaMsf+36cBNxBj18vUifczf7W7HARJHidQrlhMHZV7FvyMgjB
iiZVGSgSgAkNLao1Nq9LH61DHs6E83byOy6cUujM0Qhbsju4SlG6LQJKQfRe1NhDnPd2E8r5WuZz
hHs+jiktQFsRy/SdB/L/phCdHKxqCOGVjLIxN+K0+ps9c1ANbT4WsTe/CUt+YZ7+3fo8QdDkzIep
hDAsIonJfi571qYs73r6cipy45syAqy+XIK0BWYXdA1UTUk9HTajo92A/MFM5iWSieFUl07rfXQl
VCOsyhtVKRYhFd2aZ+INmEjySRA4vmXWMarEV3ST3g32LJ/mBWPjPhn9H354L/T1DKUfqZpkxnBi
+keMT10zVkBCsMdWnoJmg4jM5hpnu0hA6qhxaPX27jv6QEN82xcKuiaVvUQZO2/ywDZhWduZ7kYX
Tf5OtuolFoSFn8niO6aI+rQed8bg3cHqrf2VEutqfEyD7w4OOHlUKXjIDEwIb7r5LO+iGppegnIz
8ikJJ2qm7Qd2huP05gJAXYoqJ+7cWoSkG9TiEzQX11OR+hWPxltGm1j8eQMeBTI6E7tuHH1vVr+r
8kH9wcWhJJr7+rrVdkOQZBOEQBYnfa+VPQYzCTlLJuf6HKgVdFkJGujrhkkPgAHZchVdS9jSYuPh
ePzZYBZMco+WTJNWbkzX3+m3XXCH/0X+U2EHplMYP+7aV/b1F5+Wyb6mj27uk7XNDj9xWZj7NatV
dZwmpyp0Zv4AlmZl7C8LLliT5b71T7tJPvziupktjtPA8hzgXJPZPMjXhbKqYplVzf8GkB0F2Xy4
ZHyYnWO/shdnFrBdWhxI/hKsolV1wBnNOceD/5xsAJQ+eA3mzn786jEgaaWaVaMzfiNJJqhhHooi
x10GFE0Ie9qAAWa7rMeqAMpv3UBeJ8M7UkObA9zjzsLdeE/rwyukXzDrIM7Y/lnvINOPLb1AN1Ml
uxMQttF78jrHIpRdglx3UlOsNtGyIxvdS4Y3qaGfkBa40BcwvTyor+akF8S+NBkp1mL0SQdU+NC5
hBssyE9Ol8UZJOHg087nbfm/HXmxZb9jPCTHEg+oSf9jF8ZOYFdg4IusSTgql5stCKW4hMFvNe5Q
g4UX3fbvhNNL+/Qd/V0S/3v35bYSEzPfwmaFuy5+a1D09r1KgLBnyxl7vk9G9n+lVGrI+GwGBYch
Pm8ilDz3wmXWSogGODH70VQo+xYvaz8LeNo+MOFS6TgOY4SQ81vB8lrH/GAVEGNuzmScMdEU+J9V
Hfmrqn5SsKuQOZ9hgpyQAWwKNQMN1Y5Hyt4K0FuNKsMSTVIrKjNx9pW+DCL4PFP5Bl7aby8Y/4qo
HuTEf9vMtQe3mzo5ke2xus0S4O/TRKVea3TjxsLMxByL5gjMyIigY4QWxlTBubM4d9CelnIe6+nJ
QkEAduLEVErDttZd39Msuw1NHv5luR6LF65dtQFNjPAIu92g/g5iPsIWv00t11upiH7j4SvHwvYc
tkd6ShyDsdzQ+doflLyteOZrAYTFoVq/U01BXCfIrJ/j82xTKiJKzpMZvG8XnZ7n4W36+KJaBuhn
q0pkn5lJuGRfmJFBRq7XCNl97ym1X8GEbbWbVw2g3L/RB+qgS48C4XKUl2CpjiwLJyIODG3gan8/
2bE9GTyN6CLy7IuCt0ELSb1wd9zja2y4jkbV5MNLRGBPNEMIREyUCtQFi3pntYlB1s+q5BqkSdIw
XVx/Tiazzw8s8zVKCAIZrkKN5vlrs/+R2Itby23z3JJZhiZRcbWpGgIBwCzLhWhW82ekv7WOhcTM
2wchugbrcqPj5xY4SRgrHUh0JR7/Da4QlAod0d4e/RTAcvf4op+ckfzkuu7dXQpB89orq6GUELNS
d0sUHemiWjyik6kjulnRZumn/3RTLnLuEoHSGk2N/+4mKOhE8sVbSWTqLqP/xTzQElGTuFA2c7KN
Eey6eby6aPtHbmZSl7aQ0ZrdQ9+VWDz0CwoBP7NCkbWOctZRrYvvrShWkAiaLuCRLHB2Bbhs8YRp
sM/lhb/g+hnOF/rDqB3whgQpI2qtjms5rqrPtuHSppEjKjoqZeR9BhRe5CVo7+9H39ohtq5uNTMv
iCGLC97JhngNJXIDRnbFxipMOnRRMAHK/4q5gDrSHiXVAkTMDhJnsIk6lrIk82+vk4HGmOHhol5s
LblAa0X6CHirRJNjg231lj8WPsn0fh0b9khZAUP57DCz86GjYXVVcdCUlwfZB2Idsg/GBwGy4y6P
7aKwIVi+9yUU/oWgWvjPo5vTSrBwU4KNQhn4kdYh8RAmdCZRY8ONe8iUOz5JV98wuRgsa20e41tv
RbRMXVbsFhTifYfWU914//IHpOdJTVI2Vey1aPjxp7hAHFUB+srC4ozacBW35wwxy29qQ1ebbLwF
OuYpjEOTyjJiFTEYYAEhfRsOY9CPvqYxZQHpmFXukNnXVZ6/8AiLWZcTvCjqsYrp1iC+3ooMdMfM
Kk7bWJygArGswVKDsIwWS00H5LShgIGbqGML06/ycAu3fOrVfb7/f2AfJSDKkCuwaTupzUxjW3pJ
GC2MixpuhdlrCBvrk3oQNXLFulZnw221AWMJ+r6fNKgGfl6owlaGuR8D9BJl/jBYBiD07TUE95jy
cf/Sjs3TcB9qRBHIdYDORFuMRoY4Y9Up+Ihs7MLlYg4P/iDZSQPoHFUixB6rvOYeJCRjMWtCcVoJ
uGtynEHR80rIMt5m5+7Zlati7FF5Z/eVzHtqa4khXMfRd67ZLv2Iu2loMZeR6CuuKOeVsJ/Botwu
V0+wrfqDCL7aYQMd4VtUI2WXKYA6jRXaedKScXIM5bDsWTJNJpKdNyjXMp82o7QHKDWE1CcuDXFQ
qORtXMz7JcUT++H/Kcq6gux660wzU6jmm1hg4VslgPn6TVcebCCC4vs24FoB8CPuy+Tzz59v+Z2q
fGuAlo93tHrah1MfNfoI6eoDRKTm9S4p3jySpsd4RID+RtHOS22FLNQU3FCA1XhGdCMqgQhchLcs
lMsCzFTRq5Nvm13onGxekwD3yzZk76Dm52U9TqzCFQp4ZXFuUi1CGTij5yDAjdjYazCIxw2dKV8m
uypMWvrWy8OoYbxlrmglzYiGtJcTJO9az0zKgyQp9e8HKfqaaXras7B5ajepUWhSBM/rGwuBuDG0
CJu0lJ/akML1tVpF0is3/p9/kbaOk584Oj+gGeoA0iOfKd1yBOywJdfyfyebx7ncNfO/VDJ11HiM
L+uMgK6Yj/qjCGmTdkBhAAsZ5O1m5FnHmW0WWP5ldZUaMoS7HFkl9Z3qNV4ixpjWi8ZQ0nUHXFgn
WYovuc6BS9nz+nnW5NTPRNROoL63LhK4wkrrDycgIc0BXhQoAKQFfwhn7L4Dw82QtLCp7/S5tgH8
hQidm8jcWs0obWl7tnWnjqVf0igtwbala8RN7u1bYVw+Ggwv9zuMn8CDh3dvvgJLhC2IA1ZerwgJ
EwaRYBSpFYkAr0p2Z4iqpt7Sc1CQL+zxhCzzSlwZuBpHw4RViRjWRkDWWspoDPiIMTee2x52BO63
5Ca2lKtZzCgAZJQ/ITWwEADzDUPM7otmD1Tq6D3Z5YG/tvhPpaqtfd65MRVWX1xu/VJDFswOU67K
41t72RyRXb66Ih1DZGUo60zXEYfhYZcSLW9s4k7v5SDhtwi/ekIemDtsCOjnllOta5sBdJn/Q2F8
N7yxL+iO0ZuksV3v6EXtcMDfnqx56Oij7LTTS+76ulIJLevqRlnK0e/yWpTMVa0uc0uqSvzgakMr
lKkuCMNUObvzgVZC7/+mPfLhSd+lysgHyrPNj1JuYa4QVogUT5bsjx0cGp0pq8rDR6uAAhoWcq7z
LwVJscLClo8vPERUryOBQSBf0yQvm2FBSHwRl+7frxRtXIK8C4UZbFsRSL8BAEKR9GDhmnJuNh6+
62UbFCvbb5Zp+bPtG7R26hIACKE825cc64vSlX8oAD9Dn3OpDS3UqV2y6qhpu7gCSvPea7p+iQgj
/xGl5X03/RFogysJlwzRLdoobMq5CDMX3b2mI7TeQR8nmNKhKx3JWNRPqFOhjiixEzdOcqJwPfrI
SZapRcsg+uKFhHVqHpVXb4AXXN79qKzITNUw6OVz1eRc0N3510u+AUYQ7QPCi9ehmmPE3pmB4mJP
IJtGlwHKdM5Z7QAMWJcrm8XlfymR5SbmGU0AuKzX+y6XJ/IwCi5LQsvEYxkAjjlHfb1yZYAxxjpG
/xaZNzn+rF2Ufmg5DTIe/OKqAFfSA+aC6oGPuw5ZXNFf6p1m8Pb4SDk7baCNu3BTMOVdwNvEw344
P2IGSO+t4aYGDeJFHjfnK/kd6G364rtefj9Q8sXKVokarczbeaQKikD9O7fEUaLHnppBE+4uT3g9
9mfopeWOotymwm7mVcjUAgqCAzYiFlV/uCml4CvVGhWBGH39awT7999nFJVXZMIZofeO1YqBsYZi
B+M9juaUkQAbY6eBArYNl1CYW2Df4TxuZByhV0/DyMZf8v2ov2ArJZVkZji3cE6HAHRTIwDsfQNQ
IAdeT1eJfoxBLYntM7Nt3VIRHK8rexQq8KXvqgA8xuovBjGwn5ryEWIKVtFOEmaa5bcT1lgq0NhY
fgyhjz9HVHAniKPR7Z0nCEObIUglcbTwkxW1KXrQheKoYH0pm8xz8MF29CnPH3Cng5hV33BKCOuj
mLgRPR6RpDxoOWB5Qmzd7aT4Kh4u93Xfoo37k/Y0XIDB7yEgUHHeu9KvrIa9N7nzyKyjdnIuFxZb
TJO99SnXcHob3kd7Wu8lYjzk8V4b7C+Olcp/OjvX5x4Y7AgIKZxrVqDrkrMw2tT3DMzfd5o8JzOJ
1FAAEu0Lc3YvJlWkHgZDRNdXJyL5WATacQnIHgP5/Bbg98kgdcYOAXSWJVJ0MtfHCkuI/RkkYZq0
d03MIP8cJDMka7+9ET0N8hCa2xN6JQZgN/DRNCZnO0l2+F3xLmV5mhmMx6fdEIjaCeOxTKEvB1Xi
9hXwBZFswxgCSfM2aNh9UYt6mElVpoT+CTdOIj/V+TqpjkTfF463lyJD6dAD2BKVIOWE1mPqQE/a
iq2QKu2SJnyE51XStHdhysow3nYfIoiJSBNWaBLEje9nlsrgOyVIIfFpOUsjSB5qREZUb2OIz5aB
JpyqInXJKss/YSe4rGY+RlBG8DQFsXUjfoiXe+KQ8fsYlm5SrDcIN7npci0DvG03i1ULXYUhWcrV
hKYp9bKAkZkMXjkXE69OeAT9shEQg0xjJsPMpVD6K4gAT3HWudvDyx0XbsVpk05kCdzpJHyFU4Nz
AQPct07NbFzLuzYe2o8hvtWzy9y2hgrLcykfzOKsGzYVu/RuIr/EogUmp//ttSlwB5McRLT4XcT5
TOjtvTuaRbDsC3+DqWpEk7kubgZD8m0pZO7rp5tKUrgZpO2Z3xwyVEGtkBBzWG0nSMNF9/eQict4
0w8nrcU30/nRNPccYGX2+VR6zURUJUQ42S9pJhgkWLkd/q6Gj0G7Dxxlnx4IofaTIJ7w0uEwcNul
XxBA6EKViJ+76OBt9FxKFFE3PBrBRAcRXART7Bt3gsqrQlxTibMLjESLi3+JITuOpvLKb/t2VI82
d6b3UhzypWsUBtfyLNche0+yrXyFcjMVx2khC+o29nB/wvSKgykOA4A1bMgEtbwr4UTyV0ZrT9xp
daDIjqNuOa1zE/9jJ89KTBsbkDMXRMAHF55NJ3I6G4kGADCCP/iyxIKbeb2irPDYJ32KUQZ2Wp52
PeDpuB19/S48AOuytYe3rP8oHr78fy6UacqBreaUKuzv0HDhbPW+5+F6LCit+rjxGYCGCjAI1+I1
bpHB5dVp6fHhgk6NASCeisWckfG64vx+ZKd/ZqbE2o4p/H92Tm0b2sAsgODp5iFKYrpl1nOhIPnq
WtQ7d+SFbEbrDxwBkve50fEl8rq4utw+FAZwJBNig9Cp31VFvhnAL4awvqxojzHsmIYDVlCqWBKw
RD2p6Jk57Igff0OLm/IOBA2ED4w4R4lpgf115jX9wp9t4NDbwu9F44Xnh1ZIXLN8EriqeO72cnSF
8HEfQhIy62zMmlnu2457lD94O3QIsXtZbHcnmL1Nu1AH+dJE7H+ZBKcCLfEFESCpvOLL5IeRlWc/
5ZjtFabQoANNUnmVMha82HwwQdbCx9qzJ8r9jcBzHSL+Bvm7d4Y/rMVZmUnU0D4qvsWjNh+A3snb
qqTpt7kABDL1w/URvbE+FJrEucUJYvJfKfpn91KUeYOZyA8QSSu4ObuQvTPDVatsZy0hn3wRbkYD
0+yZmNQ65wiF5YVdHpNG8nmAVzcYEtughXG59xX2b5ReOyi5NhZCnKNk7gv8yUaRgCiJKM45Cw6p
WBFOm/FQC1Gwslxet0keTWU5AGifUUzRJykDbi+qJ9aol71lkE+XC1nqkSCgIFWiEpJOWbMXuqtQ
8gYdI1j/QjxAB/qx+JbDf8eFNLvSMNxfwbcH6bJ2iNDEnHmVIZYrbh2OP8gOlc1Sc62wAmuqozET
uYsOqMUvfpqBmHRL4GeZA97VGjUyljZUAVB8ecVfiyu6OasNAKl4kmL9xvr6O2oIZqfK/fq9GKJy
BVc525Pazx6QPBKIl2Q8wqTV7FjvtOFt0rPqHAo/mptLXuLuhevUWVT0go46/5mLioOCzyTq0Qg1
QmRJOXVlxd4dRYCKyINCOAQqwu9wPQeZtkeGXnbjair5wbY53wAeSzdluw7CtUtP4fgVSZM4jnNK
CRE3u4f3ZxLIueocq9GJSRMu3/3daHzq4Nqs8G1KZGUw9jfs3j6qssjDEkrDmgy17xCaRmsW2xux
ACjh4G8df3Qlm6VJJDhb1WKnXe0Ipij0vdrRfKA8P2gEJg2O+r9BG2vWRLNS54PZWe7OgkKBLTco
ZAcAC+3xXFCqzmOC57j0QYMeIlhx3B0k12aH3DHhmjbBKkLTwZzymCo2rhow8eWA7rom9i+++d1l
xaFzFU4rYIO9EESBf53Bo56mhhf6NK0u4hWVMKMNd854nMXqt6PND91TpC0MzIxKvRmOZXxamRkQ
jNnm3JUiVGy/VDoMudNPaJQLx0e5P+Y7EKzKcEeeArmrXBykVS8X5o7vWb/ZUC3hYvt9SK3Jy60R
vL3BYW9PNSAFLjpya+djkgHejyTfy4DBc9drzecd6V90w36O3La4nwI6o4STlSg+z+14EcZgoTjg
Poy1ohOfzcsxoj/kfWx87CDVSgcj9KGSj1D6AsECh1MFRRCkoDEynttEbITvXjvR6KnPpKSG4WK+
9VWUVjXLusC4wZ0OexuL0QsojQaU/ni+gLYA6MtJyO5TIHcqm6IBhjpdjcug5b0ocuGt8a2viik4
lQIbyaACcL6lezhQB+ralHgc1m4IL51B8H7WAOvIX9mznYNW/FmbtOb10llTamm2G6jpp4MXe9pK
V3QLYuAFmb/ivtSSOwTC8QSK+Xnw1tzjZtffBUbtyLB89n29OAqUW4xi6Z5+NNH6bo0oUR32p/Pf
sriuiwzRib0FUFVJav3j7qAarBL+BxhBJ5y2YWGhp2xLmn5VwjXndtd28LaTsknSE+OJ6AfXQrgl
EMaSKDA8BBqteF1mz0NpGdI0G6pmRib0vYj9uWkAhxDPJZqq10PYyDxwzfGwqoRL8/WzUEdUv49v
AILIh6q1+qqH9WpjRukHCeNA+did++ES2oAIfvTNyjlwmy+KZ93KhAtY+EvHhIMqkXERP5qANVwc
n+VzxolFY/ix83IRSh1iBfLgEmJJDlyPjrwjBOGoZDgAMNTiRO6WrL9FGCUBtT8XRK/7gCLr+0JJ
3C7bncdQIZFHISQjgy+5VfkBcTznfMwgNtmTOUvIvUMcLsofQvhf4v7y5NhMKIgVBzdwhzVMGAFg
iqCiR+EXkl/IDGfvQEFR7Vcf7pMEawaruSZ6DKTnhWCIZnqvn/pqJp4Xlen6C8I8QoPJCTg3axOq
g5vooFu1e7egrlN3kR2bOYRjbBTLfh6Makrrw/UiGCCYaKWhvTDD+fu/Hr5RJHTUAtFNuNLJ9rFE
fZjBmHBDeAX87TE/SvIKKIaG5GcB5PVWqv1ISyM+ytFdrDORYsesfKizOEPe/8Uy5PXYMycau9C6
YRgumQOBNCiL+4Vx37Ae7xxVHTie9aqJH18XFDb64V/6TP1vNi4TYe5R4uRJ3g4KJskw7YaByaHA
ygiHCKpM/tramiUE0LniQG3nLsP5QsZokShrYro9KC7FWLj+kDOtR8kWjqOJvNEbgqZoEWhCSCU+
jiqxevBlFbCAyZmeVjMQ2VPBLweMNJYMsKU2kEJbSnZlbD8cLlsOGKI9DQAppw2MNY9j1A09A9c/
R7631LBOw1mNaB1m/IsGslOzQJa8V20HRlmyq991jCo7wBAOVwEmumgNfUZTbhb6cbv0QJE0X64v
s4hLsMxqbyFrSHzMoaO77PugKY1J2dy+OkzRbtR4wGclFvsN5Mngk0bvA7f1d+bYwQgdJxbaXapR
STkLxHgz/bXqG78BKz1CNaFWY4xevjoExzZMq7ThKrDUcmPvVrjn5+gIY2hCbmBWFbgJ3FVuHfxd
Phr3tK0IJHI79E8O+wbzKtpxg/mmaDPykYHZnZcta7H92GFpKdAz/q0PSsk4MYM5UImroF3Hze6a
HI8lMY0EWVfTNlaCUWjEV5A66SE/wAJif0G/bvWkARV/iOy1rerKD85jbidnN1/QgcljRc6w0DMX
1JmPxxkn/BGRA9ZqzWzd3OUgy6ogYSvn5GYNc1RskfK9vgrBypJLmRR0tjDN6eXCkttByg3P/54M
nidPYoA6CqajE3s9ZAcbKJJ6WhLjwpDQjla5a2/+LGVfNhBZa6lHmblLpQB/jyIF85NcmMgfSHgo
gGDHNrMaiqnw/jSg26iRJl7pOcMFYUDGOhG5R9rQDAtfRzQ00ypLS7BQJei3+yhzRScOLkVs/A2E
5xk61zpbsRxe2dbpgVXQZukxxVJ1x7a5ARLjkp+vgN9sdbzAtmhmYMZEFq/uf6iN7Qcrq76NhpX7
Zcx4530HfjVS2z2QIBtAy/papVkFcAw1xQ8Z5H5TwzCajkFqo99ejfW28qf5Ka2Kh53l7jKXGvE0
+D38HfQyqWp6iGv7xESNrZ6jodpTTIZM133A9ebLyB158iFDfttKQtPXE1lirkkeCUd1GmilE2Qk
7vb18PyQHfUpFGNirnFZVnXBXS4ZPNfw12KD0xcxd6B4ObB0qWMrxq7CPv8MOb+o2EaWNR86JHYT
SDMBNjls/cfliKKwdwGnOR5ALrijSqIcwTgl04DumNE5kGkW8XRCLK1GcvyCqpy8qjeUZfWHN2km
81HydFFwP5vher99yXm2GECACOE7bQx3FYxqAmyhI9Y3Q3t/9IdadNrvWhvQ3bvc4+PoFMMjn/xb
1rgYy3EjeL90SpzhDbkt+h5aaU59yTGn0TD5sqvSSKlLMEQX6BCAbJZDI18jT+PgUdddwoU1TpeV
Avbo1+Bg5GVOAgh24Wijuu4kHne2EFw+oUTi6l4xJdyyxni4pg39EGvG0ZQLSrM4IEdeykjvTei2
/3ivVFsQ5/DNWHFVcDIOO1LqN8JIg/ry9RDVb8rGti9V2ObUz3OhuGrdDAh0WC1geXiY1JVa4kME
hmPjTI5OQMFgotvwW51eFnNZ5wQILqzwoNy6bqpb8iInkIdcAZ2W8tSGG/r7AMP0AuSAs1whMR2h
rfhY3I0ClN1QElnfgYDapylfS98fCrUcEHuK0X05l5zXWtG3i9w6tDE4NOCCw52ZrA2cBQ33xSuO
ZUzg0V22huqsRJVyKDUVtG68V4aj1NNkD/OadISlZtLEZfKD9vEJGjhd4WfXmd69NlOwm/AtGeUs
P5x7px6c5GlT3ccl4ytE6azcixRWtE7+MJa4GaQUPufmRfjuGL+IBaPONc2xHW9/n2hROsgAShmd
Ie/sP4gTALspkuOENqslHxFz3RN1dJv9WDh/ZMxQAHJTFXrQ1a3M0fBbliBWgeTXApdVtsAAR8CZ
dJhlhAiLxDHc+3IY7a6ZYBZmfaejR3pjj5QDzWZ5bTeZHNFaSQ1UtCwYdOKVLK0pBZGeZ98g9iqk
pri2HMMwzdhwtNBPukbncIdBMV0cbHroZiC2dKV+Kk6emav7RPJU3sN2v2Df3G6E9y9tc4wsx2KG
vOamVfmcsyRiEUjz7D59XGDQ7u5lNPh5y8pfOSFxbKzexQyEFTTX5gd5LowIoS5CG9JeFDJCF2df
5pP6M3CPy8iIT4jkO2KF+MamL/Kwl/MJVsrYStbjKZEB46IgS8VyJAOvLU8gE1yksIPjS77ohHnd
/5/g91p47tXNo1Fc2oygklr1MvILFn6Im6egA1rnW9Tz0TXl4dlW9l0brU532UPExem9trSWulzM
YaI/SNbE3V8FgSJm1poYeq6yMG/dGsaccB1GgxCDeh++gc43g89sX+Gb0uyUK/sWkdnzYw0FgY3D
f7YxegXZXTilkK/VsGjHPRPeidLSYpxhw0z7W2RWnaERMtmYL9u1dkHH0RM8rd0yxY2kHxvLou1A
TjoDMvSRtaQco+Ii5YUbLTW1TI+s42kDfX6wpCM29BkNf4SudKLRTHzWpBRN5Kvriv+RApNSMpT3
vQdi922xPZRkAYS6m451pJrovVnLZyY+jq4lE5P23Tzg9e9BJGI48N4i9kVF6qEwZyEY/fud0aRL
tedQV+lHeW6gAWbASlfjByM7qgKL4sItmiAzbFFpqC19Kpg8ZAhlKsJc8DttoX9QH7YULvnKDoub
EkV+dlpmsfUEPs2HflelTJifG6pE+u3nKWtSWcNQBs6qNUsXF8DgF5XSYglOnK3aovc3cU/FrsTv
nGOqTWz1Dofkav3e3vVOBNjXlIdEqBsVSpEXrxZsIDMKys5YmXW1uZ+wK5ayulMTaiJQuJKjeCYp
oc43rdWd2agwLY2qhxKrLaHAtVVqgZYaWOsU+Gsc1thNZUIbFOckc4vYW6kxQvMPYpsd+4aj9NJe
y0pYhvTJiOMwvcj5P3ijp4DAuWM/3QfcOvpKTJZXBK7NfdNGXHyYcoaEGCMZHh5g4Ap9hw4BsHfE
RXS0p9mcT38U+ouPeuePTP7XdVlzfTS+v3P9yUgMEpxa9v1uE94Hwf9wCNe4EmkTSCvb7tvH2lju
okim3zqjuqjut+IGhnsKJ35dicx2uMgQsTPzhjNhAF5pBrhHTgnn853hzbzmtWSpHhWA6q23qMhl
1KneBWndtaju2EkIdid5k7rzDY0s0WLHYr/jj0qXjcxA9aj1UjNtr6dqdDOVVfFMSOMVHYaFqlWn
HSGFXj1kd2DbZq7RMtoC28hS9yZaPs6OpZQnw3llUqG5oWyJsI80u6o2FLEOe68uQoGAZORbXD8E
eGiOvQELovX/gaPrnuRr3Wf/LlaMO+QIcL64EA8aPQKkzz/26Q4gK9ortx1qtJqkOUn3/LEAz1/H
FzeHjYdTFePDF2C/3VatnOutBZ/5OH8HCMNOnUQl25/n3/VRd4upHaOz4is9pwXECNyN4of0PcUB
/O5OyD1fLxCU0hn0pAPG/Doi3Pe0vId0M+HZ4PB6YYnjV7RCxSa93w7C/cCrI9mtRt3W/Ah7BVMO
hG5rE275KoXzqYNIa8zGdXdtffSPtqoLAcZ+Dm0UeQnpIz9vaMwlEF2NGlC3xYlnGzVe9jeSaALU
tNVvXsOY0sR0bjhfLKEBNyZJB4c/I5Hvh+x+CL1J6aLoERnTFVuM5UrS246kk7UqFe2xg+poxEYJ
u97wQfwXRY4TqhVpunzxR0LvoPWYh3aJ+aXCzfl1rXnfNsnlLLpoxEb/RezEd2f9yBZguB+74SAr
qyu6FnHJoburR1gFDbwBjrJLL2kE6IhoHDR0ZkU+H2econIuMtN92XahbowkU+QSgJzaFS3/mIJc
fIlqipc26jLwKMbNrdTtCjl7AQc0srD3Qdo5tG8GScldh+P0ikv2mPVCqMA80oLQTJk4k3SE/APb
iQUVsNGCpOoc8gSaN4ZZDVSF5owt2BXzSDnrU67HFljWPMKrtkZf0UdKN0JicIG7oO1VpexbagVv
NwXf0g4XGed1SfQfwp26CsV5WCrVFvhNIvJn/p1dCDKY5Dt5WvKWAf3+4+DOL7KpSIfJAlFQd+Ky
mPhEtJUSUKq+CvoQI7mhNlbUyZCHOTHafGh74LMN4sHa0oz7FwYB9TkGv9yoJaTMDmiE7h/me+UX
7oyPWxQ4j6NhtwefT/nKhr/WNixr+XeQdXhIwa2VK5TZ6Ivt2wB9ouGSI/0jMnxwVTJckm5/J/V+
iUQC2aaCdX024H71z9egpbsuzZivKAypjjN5xIohR7NEApT1XCzW2iN4Jl6Q66BY+dgku/Hbx8Id
PeNCh0M6YqYbYt8763yfItRAoe8n44YW+wTnLUX2u/YoSd3+kpMBc76zKsMxHqJFNJu8dn52suKn
2lr/bbPqBO5iVYQfJgnwNc2YNIkM0UCKI+XIue8MAqEnANBuiggFGQkAyPUpEzDt0BIch5yIX+ay
j42mDM4jK+h8u+ocd8A5G6RIxZH/KBuCFSkMTsuI5e8Ak7qdOYaBsgi19xkNExrTjv1Ym/323dVx
NgHj/FrQXfzngmUTOnVzsgeOcH00mgROegqnVbz0diR8focwN/vfLWUFu66rVSYp45s6ZQ4ahaeV
YLrJC0Pu2qaLHz/PMCYr35G0QrytOoYugRzgRRxz8O1nH3peHE7g1kV2DGRPvpdejSXsqLOiFWwS
42PV0jm2u8Lfs9VzBcCSF0947VJ6YuYTZiJEWP2GVsa1VwVNZmK/VEJbALVBU5PlYbhSoL/5Gc4l
Ptcl1jaDLCWmc25qIWNvX5Xjf9j66xjSXGfpyOFoOo7X4iTpIW2KAk3sDlsXcRfGOl0didnEfntN
liZI+EQIYrBxacdIhFtv+yo2/XU9XDDbGkA/X3rjCTaBMb9ot2B07R4Hvr5Hmi3vbuJp6nhLjjEY
HIpXDpI9N0pC6xHK/La6d1dhUKV3Im7B/0tVT6+TcZlYTwUbbv0C7PLoinIJEpU8q6bfyWjIpPPk
hj+iQ/OcvNvTVdzEGzTFOP/IV3cBj1hwWn96OZ7PXe/wF6zMeta30hXrNGDFOb/J0K4Rf5FJmajC
i6Sy0UcgLDwuQ4BjURtBcBWlNSF1+L/iukc2SEV5IxJ5M6GpGmy1NAKvudVZ+nuGk1kB7SghsrgM
mnHYz8Pf0mUMR6RpKhLLO3l/MXV5/Ol7Q5fLRBR6sU4T59Vkd9pYMlL2tCgAdBpDF3Y2z0OR0pBg
8+x3ayo5j80q4Rw878cHRZJ2fmHJVnoc7do6BI6mIscH1+r3uNEyb6ADb7hgVlg5j0+k7blIl17V
7TKtKRA/Wn0EcFug8irMdXM9mz9Z3m+Xlsr+/ZzrxadROPSJ5b2pgTQUkPqrL6bmQjjPoKH26Qhc
hQC2RygmBq9zEJy69imrIY700kaUEGiyIIvzgZXLNarDM5a6IixF6RckxvI5XVDyvnc40fzpY9Bh
bqBtALidn2kT+gjWcOJKdXefxMKYWceZuZnvDer2st9zD44E2lC5dK2pKeqAikqzQZ62l8iMZNCN
j3WHcOUEjuHKZfyWtiavoeX+27DcR5TwmRVgOvbyLgq/fPjMjGj1gXiRpY/oMlpjpUFJzzVfGYdP
ON7MY4M7D3DLyhP0A/xRz5N3MrbGRcB2P28Wt31qV6kAZVnPYIRr1x4emmkU9GR3qoBCaE8O1Cmb
N+DO6CzbmIY5/nqj4p6EOvMnpgZNstQ12WAoEMl49qw2YbmC0Ia4pPEIbIsib4hE1dozI7hMrdcL
6lO6YAAerwFhuFGxqB0AadyaxkJX32Jat5Mpm7n3lD1eCRsBKiiFpTyRxiRM3Wzp0pN+E+DF0BKM
rzbmKhvpaS419oAcE5sEH26NQ3NkwsfD1ZabW7A+hOGq2x9DWwy+WNkhsGjP0quMLhehnWc2wPtv
Itxtagg+zbyHMLtvF7hQp5uUbqzxGFSpFD3rQEUORnPs/b0BV+IYBz5jYCIFUtW/S85yiKcFp2Um
Wp7YGqguHOX5Z04RdAQyea4kCABnmZMY/aGH2s73UWRHI6kYrxkgOcee+UWUVtX/KNl1iQKyxHfm
NYNBn9WlRGA+RqrcMSqt4H8/vBgvaK15lRcRmeGcdvJiNPrWE+22za88zl+HQSfTW9hhGctDlHUe
GIxGIWcRAv3E/TNftVUOVKSJQRuiIHD0LIVsxO3Db+tNMQr6mBt8oRQ4t8AqZOAA6tEels/CnNGV
meGBJG0ZOq+o6TBZSp8NyDLSQRCp8ZTyuoCD6AXq3hFQQHsFnlnI2GSNzqkbk83FnMXIWE+uEB3U
IuHlNpdzL0NaqBCMj2KThET8Ye+nxRFGY34XVuFLhm9/7qL1R/2PZdS/4n3NRA0mJaqah/cCDkj9
iXTCQg46nmUgNxh0Fbz/4eUgmtYObFgj8pbACKvZU+AtqWmpI5CrVleaJgdXUMq+PabRS+d06103
eg5CwgXwsM10fVGL4lMQGrF9osKBlhnhyHToSQgkPaS2Z/Yc2vwCcTMHg8drWU2Iihw4c9fVJqcP
wc5EceRgHs5FLBmPD0DMeUrc53aHv2N9/QVm5yQ4dGJ3s7SNeqUPd1aweRY42MzwyIdzieldQVGL
+3Hxy8/fpFX4NnqYsRVgL2CFhxDrDACpfcTffzKmi6jL0AiSzLVJanaRzpjveztYCgLcU7NbhPuz
5GBmdb0ggNK8D9rqgKVuFxSE3R/SK9suib0dtPwXLabk1kyrDJeDJo8dw0Pgy4w+hpQLMyJ4vL1c
PvE4uCk8TqpdCa3JQ3b80lWCD5qjd3jPBR06794/xzWay5VAA0OUJMgfdpK3bLtiQ3NR7ZSb83Rj
Yu6L5n8zhBO5mPX2q7cbVHvI5Y5eX8aD6si7VuQCgubJ5/o4t7NmyuwXSDz13u3khfWKrQbYm5v/
Kjf4nyFahK27nolWssg1i+Qjlyi5+KYP7W5onnJPARk8xsiyetixWXmwHV0yMls7LAgz/AdQIkmM
CLnGc2YDeI69JQ8fFsbeF0oOqGwr1INV47ROnJQC6q1FRsgSTEYzPxRHQ3DJjv34JRln5bvHps6X
Cp47qaJCdDqPOpzKB7ceoMD9Nihn3JoDhHD+laV+qpicCHeBstII/qfe3cvbNPW2OXQcrGwo924s
D9gl2ExNdpqf9afusEovwvzIAjS3scuUM4jKRWAczbobOswzGJ+qn01d/X9LxIQSJZo+h6/fDZCK
1+vAIhwUUTijqQk/mmIqrv9cZwchJ0jdI+ROD7Nxs7EKpITzjKgQd+1vVkfo+JNZTfBa+8mE0BoM
VN6uPNmvwGQNBBCAB81BXFPBXPPHrAjxi4xY1OYGoymwglMvOAmbXL8wjir+OdWVj5k4TuxdRaqr
p4bUsEbfvCKKt/MrGA5v05ZuG95VYAmlNTRGo87EMu5YKp8lPGi+OhDauqHodHk53Fpwrda1+1mt
1LTQbd5eyFdGmpwZt9EKHR/iBzZPyKN31G2S/2H4yUKMwmayUPbnVplcDEZYm1qYNQbcrfiORPRc
xWoCQMrKFsp6aZBC9tpLA9z51pnsBFjQZYOAO6GCgbLoPmQsLLpT2qgP4mysqeSpCokU8FokLyJI
VwE/sN7988Waj/J78828lAxY9lfLBCFq8h+memmCBWjs8Ssyo2WNDqJ0Zh3Gz2Mtx1lWcX8q0QCF
vb3InaM90gdcw2jTk7x8mIKBZiw+W479vjEcXCR15+Nyq4Fl+RbFVuF4cznWTlSmPKIRHOpSR8q5
cxPWSNqr1pbV7trLc8sPF4Z4Qfjb9zTDp9b7gLeGOgqam0GXRchUw1RwC/i2dRzc/wYJofnEsSh3
JzqINr0/wRNpdy/HbnmmLPjLTbTd+WuAWkD4Wr61wUBrejlOu/8J/Me8/BGpWurv0ZRKnT/Gm7Rk
6S0epKmeve5SEzkp6p4ApekHJDIz+2ZnQ6aAePB94QYQRaJR4TfY3dD5ZkD9oZeycH1Y9GQ3QIEL
CLQ2dNZUiGKEexAUiq39JHogjcGV/s5Jepx2BVsAeG6kDaf8FdIZspnbZaNTai4BhiG89T1K5bn3
Y76ipMgKsFUX16xhzlZ6d/GESEokyeU8EckAgdkd6CMFfq+IHsS+MSA54b+JwILScauFgAfXCPsW
jjTRmZ2fgltxtg/YoYkMx/SAHA4GXcvT3a7nVvOhTod66ZEMc4decUDsMUH9JCwa1I7TNnMi6yCp
VHvh14mvt2vBvaydVFOA6UNTV49CRsCSuXIWGK3z3Phwa1i+l6oeqxmBcf7c/1AD0b3bIRwwkj9z
p4S/VCTebVox2MaDqD/MnawWS8ldTCQCW37SNeziryLVBnhZCaNX6EW4i3s9cjgeAiHjZF3Kydrc
6HLGiRD1cqU14469++9Sd8F+MVjwDru3qmZd9LlNQWf4Ze/WBGb3fdPXmW23Bc8kZVOnOHOTNx7R
hW5w94z7ukYI/CyauNewHuGwx/Wvrnbi8WhgfIm3ffNd2RucJt605GWga6d7kFEgUhsNt69RJHf4
Q+lGD1+pqfTHlFaLWBFhfh8ltFHjBSsOIAfGxJHGVKaDlKvI/D2bTb7wYfABB37u3X51WLLdTHya
wJGM3Vv1orYHZ2Cx/RjotWkn7bLLdSG3YiZ/oI1/ErOn2qj3V7ElHHKManSftqvvnDFylNSnyePA
X81Pxr66XTxwcgIpggEcSfkkgdIeZvuqeVq3KFrAY+ZI48PWW7TTbF3wfWICPswA+5zGNYlrC5Qc
zRkn6eraDcthWIBspMH9tTBYmmSzy30ZS1dvtovfByOsHvO8IkGf1/979VtQtvpbUFM2w+vMi/gc
0BeTBDUQfO2imUaIryZnSHBwX7NI+Ed2ExDGgKO3Q63Rr8nSRBcPvaROdRJmkC3cCf8tj6RIh1gV
HVKlYapP9j17kkU80OCYeBDiXrwESYh8RES/O3wVYm7tTTzE5mZx769CfSQ/HrCNxrfBrLUnslOs
pZbEMPbmXIjON+7/hQm7RvSAxmGwh531U9S96jJO3F0GoNiE1SJi3/G8wwoFiFpdtB4fI579JwZV
sSLylevuXQK3Kug1pPGMYZ7CwaYFIy/W8lgYvMEudxTDpU1gloAZYTHS8GSX+MMpaZX8I0oPh7jf
ZnrXL3laWE61Ou1bpEujunIBlNq4wf4NbKxr+aA5/a/tbALL9MLRewj7WJtbgX9cn8jn5JRser1h
IRohag2n1KdWK/DUW16tXMXqoGZtOJmqPkskSsNUbEAfmDXYFlnnLVhCJWydPoXSBSyGrKB2HUkA
yIMrWi0Uizn7e4dE6HdBJIMq6RS9xPGR9LbAppwECM2RekxyoLw5KZQOZs9fy5Y3HKWg0iNilgzi
zGhUL8BTJUpQkXDGdu+PiPqGIlgjARI3qOdhMKHGzIn+ACUuyWE781JDMr+1SJMHrYEFMnHsvnOt
RDn5sWzCaOEWH6q7b8uWyhHzYKUwo1zqkvlousZh9tuO6OCWBDuGUp7JLwCVfRFrNrZJWDZ8UH8c
V7QrqVlsDVs/SzudSzWYMrAs1U/b94wKontcMLtW1dCTmroAnECNGJ3zNm7CcOg1r2MKI7T/xkir
JweFJ6w5ra7Ra64SJYXb6Z3FW+Y1O1CbVOWdhbA95b8/rwdYZCX1QyqZ0Aywv1AnP1I7MuhBFrNr
75/ljBCkfUls8jKobmK9IznvU1iqnIYxOksAjGk3dGrw0PCmOMqaHt2ml9kDvtQpTzqzdIs+uAYs
DMVtb3Eimoli9SRkNQ40rb+4DNQelGyzEpu50r7oT7rDijrzYZk3Miyq6QEMKqVXL+7GGCYjc7ST
oCXc3zfij5jXvXe7IwwkwP/emSWaRf3W6v5u//lCHartxpTCzaQkq5o5/BP2g3HJPL3O5iW+C8fB
V+LxvvCI5psjKm6frrBqiLsBuleRRKKy13Y/xAnmCD/82ikDcYDIBz+JnaFvyWq1QbifjEQLUE6R
DrV6rLM84U7SaWe5dRN0XW0D05Fyu4wHmGS84pX4GwTvsBwrNWhTmKGxv8ZoUJbaLHjdWLdzNYnM
jjbvcl6Go5DR1jUh1RQ/bJgx7j3ayJGW8m4Vz/TZTqSkvcE6MJiP5bfnLVvb9FV9JEpyY1Q3TNBd
DOdLiTWYb8Mya5EE6f2ZCFzBaxelb7DXbk14pgVx9oIpPWBibz7YDtXa1j0Ru5h9i7JYolUwV9Dk
5tkY6+3u8QtmRL+6FYsXCM97kEIeQEvqlPj/RTvSIL96jREBMj7SfJLoLk0QGp3ohoJOL8zJMa7T
eNLKvc/Q4Hg2yp5YM38fpO4X6pmZRomztqlbdu2EGEslY2GwyHEc1yXDEvUCDfdLurLdF+pDzagl
7NUlLgA2/trzlbIJOCXfOiwC0pjX4P7mReSKE2QclfvJgSX/RxXIwodo2YI+5mE1ZMQ4f61Y7ijS
v9QaCy7V6KUATBLTu6B1bUDQ20YwydyLkUAPTNuOgtJE3WSpndreWdjhVemwlEWx9CE7q/oZAgnh
0MXtSjLOgUWBy3NqHJB/tNrH+eSsdzUpkXjgkWtdQGKSsC6QPDvKPIFBS4ydyioUBeL1LzSgekb5
TTA48IijqOWW+k0TCIIbzw2l1XWkdZsyCQkFo0p3cz1j3DGDwmWa8iD1W+Q37/qKhTJ1Ox+AHO+5
CA756kV2F1+PH2JsPnj814cOiPk8EE5YnHdANyqovZkZyZrH5v+Qvsp9TyLEnP3BjbNHkk731XWZ
4uyjGGsBh4/Md85BM3GyMygBLGEMxWBOMIwfXW8PZ8bUDfUduG52tUr1hu0GRTkLD6LJ5dr28l1r
yE/Fxf0S8Ej5iNiIkAexBy4VtfabFKselpV7hkvSvTZEWLZgDCH+MDaqhDAJynUI1eM5UyrZALpM
Kq5kdFmwQYenRKnXO7hXcusr7DdfWqbRnOXI88WtxZBW+3b+OJPf3+/awPU4B1xcabBA61otHBjK
G6p7DOqMSgHVg9iV75NPO3pqCXE2Hdi7B/KZulWNKOWK2Z+Vt6zPxCvJ3HfEguAAZgUC99PoUbs0
fFU2f3vX8ZpVLqnCf1II4afe1hoi/HSBeAz/bmJcxARb97/tkhxoUL42ZsA54lyH7+XOTVokFaf3
LAXvkwywr+ahLOumW7QRDVP1iCzP8MhXwyO26NCJ7FaSucK7Btprd5+dcFaiKysZ73zqQTnFUOKZ
O47D8FMfun9M3Eyr19SGLAfpM6P2sjApFlTI5mW36vTFa/iYX5/9JGbee4Qg0QSUuaOvrPnsUd0x
4MW3oKnwlu3RyCDbwPdplLQxuPMZ1sLr38bIgl/Cz9t16VJubVOpQMwhAsVltO8z1jxPc89SN5XI
esT3y5+2Z9EYYInKHY50YxdyEaBuf3xO8wEmnDqZjCZZ0WwDgsNpxMB3eE9kwJmD7+QR+pedEDxW
K8k9S0wmOen6olLguYigx7W3rx8qDgq9k1C1Wui5ObgXcFlxaD0Mz9C4hiUlazP/fdPjXY1G+3Ku
jnidnMdezlyzGsNuoiIE0HigmSVqucgvAVphSoEbgaosLH1wMULCMcWRyqQW7tqo/v/foFIwR5x5
Gbf/2uSEs3jFA5fec1tBXwijYSznQvBvzhmf5f3cgBL4+O4nTAQN0/MKPXZFIhOyED1C9+YyZwvj
GjGkM5fP1T/5JdChRAbprwMzHShEsL8EYTjRUnpM74we0iyju1IKSLOWzk3Wql+oYrsyrRXbVjNT
jt1m8oOSUQcJXMW/rCE0gCNZvCqeHfAHc5WXilBVzvE6N9DEW3ZsxJwbe9Bl3xvOkx3yFrgvcCKP
mJ2WaCST4yWvSwWYbgEsdzt8Fbimz1TdwGLXKej6UL8xruSZbmg9XP8UU28Jw6f3hMGSUDEEHAvp
aC0KjocMNiaJJKQw1ytAJOwjMcRQovHd/RMH49NdLzj1E+r4WfRaVvpPvAnKcN28xkJIzUi4Fcct
PTMfXg55+NvCHJH9BJz2WXJBlYJDRIqlPg1HQdsA05GtL9XCJR0qu/R+EizzI9yGg3tjLUjkVPYu
pF6vDxx1EmOIFPkq7I3JfYtGngqqVwVvNN9Sc+8osJhCAzC2VtiQGWksZQQWAG8xRiDxzAcANYFG
VFL/P7gWt+be2x6qJNagbVqdfN9MAXuKHlHeG/DdkJx9CeQUP7W9pQkG/S2Tq+PX8AArysy9DP2N
MW20FanUMyoCwCxmzFGFkE/KZFM8FGgRzKqdiTovvXuL1nZynL/DyWSXVub77qkLB6EQmjO98rDl
uzMNbPE0/83OPNPg8Q8ZkIPyIAFRVdA14ZJwU3xH//F6edhqeFK3ozDawcU9p+dT7fQ0ua56aGP6
DuuZdTdOKqdjIUmU0BINDp8v/CAObgaEx+wQGV84t4vfmxnFxKgScKFVe83zYqte8ecin6q78dLc
XXnotKAKm847wBfumuyCDNRvyo/Kfh0vwfx4L0nlI1DjfuH0HnzrHihrkGMjaQSMy98l0j6ZP0nG
ORQDtuHNGB500LDD/LQF66wrQ058kMgPqaW7mcOBlFFwhmF8nZPDt3x7+c68BgKUJXqL/bonH8+W
fkjU3HWzEOwb+Sl8iZ+V4FmUP+gUD4cWXtNTZhtL5MS525fQD35zz6YPHnC+l+5FYkZuJOfnaSHb
/Q7hAKwvl8mobPSr9MHzzVGTV5Wza/DtxgujkhUiw3AlgRL0zj+bbWR3BrZY3y2zOB5jCq2xYO5N
D6Zw8CGYKVx3zsNyWunkihnJPGEaqY9L817ea8MdZbSt+kUX4cZji5JxfpHGJnzWEy+mE2UU3Oqx
ZVR3w1dlbL6sE0tOghgSmfxnNcf3oTHa5aNoIGzEW599DyYZNuORS+G8NzMmI/V29WzIVOx2tk4b
F6vK5PkPx3rAUPNs1RjqioFsS+JuErLdx1wQpfWR3Sm0xtMn2iZSSUjs8ECDxk5G2HhOxEcb3E1M
WUSmeFSDWMEO68027KYF9+qqSRgwugt6KUUidqLCYUfTpLuZgO6SIkYWwB/ov9ApwpaJnMtcCPOQ
NRv4ZLdp2HUwmpjCr/c7wubR+KhDvnGP2KmNxxgmh1tIySdlsps8TbeHM65H/HCepvNuiMyG/0pv
r64E9AO7tctqes1sECTsEo/5QmqGj9fsJeRD4fsvOR6waNps077ax2mYzj0MOK3lZ0/7rl4Gapru
HRgUpA/lSH0VVyrTxZrKPWqWOwNCCgHBb6uxfYW1jXi9m6jxvd3hXRRA23ZUV3yOO2H6GZ4qIhR9
rXVjy11h57/ZZSCwbLtolow4YA69td4hBdASm8U9kpMFJlpust5xFRAqzTbf4Ny72fH5Y9O5GGmM
9S+omOo6yoCoVi+e8qLTIr8KkNlneKuYoxu5dKQlwlFLRO4AyTVX1jrmk+PW6P18PwUuqI3WicB7
b7wi/0WphEaQPz2BoSRQ3Bv0vinlH9NNKHd3YVUSQVh9CDiI444Igwuvo4XVIAwtqg0cMpY9zUIS
70b59LIe/7Bf9wUrmJW/8fxdvigcqiaV+sdYx5M/r3Rjd70xiZJvceyfKBvDVKdpSkPUvAV+HXv5
TDs6zIgaD38MObp918yGX8GcKz7I2+7CLbxK5pq88gk93TnylXusZ5RtYiiMEJWoum4E8nOy/oeM
rRbrLSq7Q6I5Y6m22fusqAoS3SGaz5CUwwIJ30R2EW0YNtvPBeEcg/9LKvrnIF3YExK7+QzgfgaB
5RAw5tuSKRkZhP/XxnAfqBYWtdwbISnYhBQUsjiGr0Q19im4nYVdzhXb25UFN3ADHsSHh9PqYcZA
aN1GpS07PUKWHoBnU7hGFmVdihE0a+D/mBtzWYYN8b7CuoOxIKCv+5ROIysEhy3BFmKUiYvCs53n
KW9Wj9INyu0pl+z4MvpbTzuuZDTmASkHj+Uf9GFBJvnY5IETTu4BHoLy92XOHtFVh76ujbUcVfyu
DQt6K7u28M35HUWXTNSeiYvacDiYdAv3yPLHTYV+fM3lCkWGsRpWu4TS7yJObfvv3CzHsLn+/NoO
vplynl0QCQJob3mK99MRp0PFaLdmNufNuasYPP3jL6626rxYxOnbrZLpRWGNLCNaZIOE6Pcnycr3
hmwhhXWt+fjQHvmFzxmrOUVlmzycTwluPU9zA+DtNiP+zb9fl2A0Ox8UpH2n9Dzm5ajl9ar3TB8J
M0CmtWOcCi5mBgIzFnbd2XPkD7cnGfAkV67Sid9Q+86mJl1d9rCZV7HmViaGX6TRcUpwoXOEjocN
lxtkAVYwfwls16QJLPK5EU9ULRDz0UeDTwvaSYLEjvDqcq0Z1WW/Xh/fbtkDZ3NLCsr+REYMqqPn
NFpSgAQChxUrWaVRiJMtii60E+FrxlkJ/NcF0ocO7luxpNyOdRpA+ZbuI0kiMfAADAXelQs/pmJT
zVdrUGAEPxZmQYympUxc6FTp7yBftao9Jh/4hNkXItOv0pjD6BpNWv5XIU+Gksgotxet8oi5csb+
Q/I31M5i8vZ3E//4QSNmVRTdps2bdSX+4OXRMNTyeWnvZQoiRjEzkly+xdNHZUTsXNKt2Bqn5yDk
2JIe2IvmBTRwPCdy9uaC1p6NDbXT4+zD6LKkIayyg5epyELfC/v2drib+/SGnPQGUcJJi1uM1Xbj
jVRJ32o7jicy987ZrFWxr/V9Qa5sy2eIaSZEs7gOrY0jWGmPtPMMSQwgnDrw/mQ8Vg6090Hp/Qnn
eWFPTzurEbIiJxPzDRggyE/sMVh4hMj2WOBzOx7pT50bwM/Ere7CIPPgteHDni6hlHlmrvyGivnc
LjwyXib8Sv7LOS0VQ3TKXQpedbm18UFvQSOWjV2plqQDdvk6bvVfTTGPbUnOrSDBIHXErpklKLby
EICeqi+jE9P9I/3CkF+k4MA7M3JSingxAWx+lb3jz1S0Fu4jKIVzFx2ATlAcidO2HZieorbXdkqB
tupwL6+SS0WN6d8B5p6nlO+GVNIKdMMyJU7seUa7Jiwx95tUwVGhT9lvKLXICohZvtRte5dTRRI/
HfLTZDuzwKfqH6chKtlZwlCtOTqFINzuLt28R0GvXo6s5c+asbfaQGYqsF1lz43tMqGCIhTJNUgh
v0AR36Fv3JN2lGbPDEcdyuxHSCP8zh+esAOuYwW6RDUTY938QX31Q3TWH6/khWbEUpYZ3jcMnSEq
K2TbhZ9iRvDRhyUllCZp87zgt3GIUEo3by8BQthJz9HASfO5AClmOAPgGZsglCK2H8GuMufVxQFX
JRFjjBAWfz0g8Mx3sAdxRH4aJeVJcaGXbUztVJps3rgplg2mIXSrC/Vo33fCE8QiI68KURhj927S
Q4Ws9vRCr48ZFap85+MShYGcofKBnr2CVDj+QdtvuMfQ2ISlfLSwnyxaXdKiYYRJGpzlgcxbB5aD
FPMvPbuyLXb2fe8zewdvUnSubLbBt3b3AMFTgJaz0DzIguJXRBTPAsxYCT/8Uq/lVtjABj/cAO6P
gO4j3iRydtmyAJYQLRRTPYjwyBbsHoHxBr5pD+gkGg2pVv81mVdjM2RHguaoFjlWUTsR3t79J560
a8Ih2eTMsZ9gA/TArG9n7H3WXS615s/oiVEO9p4/yH5uZJVajnlnFchKoQvTd4rvV+1dNw3BDWUA
agf7gW+KazJUr2E+SEbjrBNcDjHhfnF3wryCJFJFnluhr44RCW5MsA+zmwR+YwgZ8VVFDvwRlMPA
5daMfq4JQYuGVjdM8m6tVxCbR3uRagLnvjZoJCQofakxEVOynxjWLwVj388fCqdStRnafFovO+F6
F8Iy88Ca+DR4pICPD/4Fq/7qrG5vDQ9YryiQq7ybpMSk8nyafOcNqYtwvlXHxQRaO+81/eozrUMa
tK/fOcVKSGE6zBrbCrezyomNESjXmTH5w8CC83mFypP0Gf9m3ng4b9wmN/BFBc/c/Ak0jSTefGOl
p5lZJhtttL0zoRZeYWiBypcpPbeBSHGQAU98CkF53KIHQbmmcodXwZ+O+HuzxHNfHaK9LYqG/Lt7
PSKkQir12uoNli9pbu6P442+GBRW0ENLCzI10yp2t8y7VXo6QFUA91E42Tk+q4KgeiSCSrJOd+0H
Mqx52JMcDlCFgCj4L+cpetcxBEo1HjwUxQ252DDYfbX+3t3hUSWpQyttl28Vc7DPISKK/ahR+bny
I12bz639y0WN1U+Vkyx3dTK5WGHkq2PLE8Rpk9/wwFL3rjhLWLY3gXfQClpdWpcQUjmrKCvy6tzA
c7mdF7RhpNV4RW0VoAEF+pG65iJgWbXhsKgc7BfuvKmGMQH4WKSKpMbhKl073cPgt3S6SO7+ao8w
OtulxyT9QSdkd+XF9biqtX8yV3Jwwx+3ggAVRKm6b6BWHOQOQUmoSuPd+hL0LV0hUwiAeUcWbGap
jYPR5/RDF97BvISzRhmiPcbr9L3mY8dgFODO8ur/savp+u7w8Qn+2QKMeQhFm2xju7zeyCUeXDTz
HNKprQehNOrz9BQo+pyf2DK7MGgjawUPnvphLJHyxPfgoK+EUPPmCIFRL/4uxmy250Y5+2afXnxx
K1Jtutu1051ccffPogGPQDg0TIMjSnxYY8dd/lkoW+4/XvPryOBEq6X41gKi426oXvG3ef+aRZoA
9xXBhJ32wnSOcx4hfkL/QktsxVIjMooAjLcn3IUJe2Yj0GCw4np/IVNfubRTI15HSTmDQpKoTyQX
MyStLDZWsV7SLS3AWxJ3dwLHH7E7mPo/HAWdNQ7Gx2CemqRL58pUMhtGbPJJGd43pO0zO65CKvo/
MjcKVKkziUkktJMU5XcymkW2p2/PL+ImY94KJfqwigc+Ir7+XPs6IRvQniPflFfAsZmWXCzljRnN
79i8dNp+J1RJfqBOQR1wTHHb77kvd/VLOPlsLSjii/81al7rpTPbDB2HOfdmOtAfJHxX5QWMU8Ai
nUZNN/ZCEvuTBWKM6C3m148iBlFu6f0R5FkWWZRcpah7sfJ+Hg/YSquWHHT7ClfSPd5iuVmTTEIP
68USDuK+xm/NkZFx/BxGPcp6ORl8kgur4TEGFoeYnoVxevhjMcsVotxvcZqHl7oGZ8BqazNUFdRQ
aT/rzTw9cuRwib/ZheFOaok2JbPTrhk60ni+15BI/3hF1GgaznpcJaQl30ESUhdrkNzEu+DmRnHb
Cm0ixBfkpeu2HiLlCNqm5woXEDxU9Hmeoivv6zWd/aeHjI6lEtI/kw0lGYgNe0uPw9hvnTKaQX6n
ejf2m2yeXH/9Kzuk9V0z7RddFXRI3R0gNma5qLRBuA4hu0BOLq98ff8fv9wjgDFfU77IqfYFKt/F
dR03vNveCP6JVd8yKJdoZeeXX+PlJUlACIiBmj3XDgsPb4AIxou/idtVIY/ElQ3KUV1tddHbt2ZM
s7QKpBO7nB0p4g1ZUvOtr6nTSk5eW0crVB0d/GhJriIQpkndJifN5H32KjlCci0k07mGcozmSsjC
OYQ3ItbuYlU7HRMkt3jf8t5OhGPgpX2UkUF5u4IbzWLllhDqV457s5DHbHtkWvjyuP0mDET79Aal
zWBaYMnBes+l/tgn1ueX7Zk0KhDatGDjCm9zl7l3WndDNfQW6KqrfrqmBCw/NjnNmjDg6mQ9W3xd
sJVFcjwMouI8jsAP+8kNwy/hFho7d8Y6oVn77lQjkzfZlHffY6VFNioSd8WoDkqlgMAApGlzbE/Z
kPZAY2gcE0f3opDxju8GVC1DUZgXgn03/egy5611t3vMZ0mYjbs9iJ+8Xx/tW2AMfyespQ/Z1kRq
LMntfGoGVfcqvG8lsFfonRgYMa39qqFTIIrbec0Upxi7legSDweJZapQNEiJtsZZN8so/qEZZjSJ
TQejParXDC9Tlh5cLaSwv5AC0SOKfWxo0ko91LPkHhhQ5lZZ8zI5Mqi95pe3bolyHcTH22gLTOwW
Og4TzllKMQiX3IFnXD2sO2Aco3Rdl/X0YjjtMqP2G0AaNMJCtBLKYgvZulHUk3Sq+QeCajT8iVt8
GdQT2Dxlf8P1b+JXHgpaUsJcM7MDGPGHcl/J6OFDVcUZCRCgmv+0aSvi0Uoxumc25zipnVhFcVZ0
2aFQnOeilo0m7i1ETcE2rJv2BLMsii+3tlIjKWrrrW4lOIkKicX7BdA/p7ArhTZi5/sVpPg7tj1Y
8zw/AtRbSE7KAWn3gCiS6iJPykpSd1FdX+wyl9kKc93BlxHavKf7ofn6mvsN0OHweJkgDjRrCiZo
fHOi56fHafYFx61JNCvhGqN6K/sBC4otnaoHrdSiJ7qt0HBr7Nbdh990wosea+NPtKeJ83zMukc8
ck/qMIJe6Hk8+AvwyuAtR7S0urYWz3TVW7eNZGYYzLh0/WjleDWwqqHkZyVO+H6aDXuVo2HR4SgW
2+9OMvRyy5OdyVR9109qrM56ifOo1OlSrpzp8L5nycS21TABncZy/7RZ3eB5p4KNlGyj4AMF1pKn
Y8QjdiOzJ26PBK2ht4OS50bv/mZele25q//WWO+1wz3TkXCqLSEXt1E4klJ5OoGnnEQnqopMZiSV
bJbqIT1wGGKVEVUTFn6mgFTsvRfRzxim0gGCweHpPB4+uye6j8sR6zpwcWV5DkaJSZ7m152r9c2V
S+8UTzQ8g/LX8fK1FEzzgPYMQwJCqaLdNv005t29C8HhNbEFLL1FgC7IU7xIhAOZ84z9hoAK2laJ
iyDpp4ZJcZYfz5MshWB1iZ9PfSPROHrixmd1yfM06+113HJY5YT5YUcIPf7RkH3d4VBf4DaFFM4O
efve8B1yuG/2UrkF6FixaeEPAjanRJPRtQULF6yZex1gbW5YzeJ1ahTsv9PL6F2dfDlMDTCXGyNB
LuUMj9o0+uFO1dnfPr3Ut9jVJDrKjCkv20vtIkV7+mdmVJ/BfjoxNPK0qFjbKQEWMwXH/d2pEDy0
UYyT6IRkGbRdWo4MQ5unb3HYcOccl8yoFR0knHAiKshOXwjxeqCe3QUvMoZz0Gio1+GZZex4wAYX
iKWEDTRBEp3FsLIzh9ZS44Ndntee+4mOvchfEpUjsbUBg/eZX2jjXqRB0jyf8iQT8rFW8yuGgMkK
vxTiYeSyG1kwROdjfNp1+74HdP5PkR0+pG8TtZFwjQio/HPlQrXhaE66u4c1OKIRlymtoQufJERa
pXL9NRl5P2r1VLQO50if4vv/x2w9eW2eqf0ubXT6wPHedFPIZtlq4A3JwOenyggAHT7RYQY4Rncv
5mzt470Gqn0c42G16et7whYbdKDvbSBFPDMCnnM6fXCRhweAdbg+oPtJ9Koi+CMN9GFOW5CYGvSK
qSnv5j/Ewbhw9V7pXjl7W4Xvuq2+ueS8ThNY1pPvLTmoe4BNhfHtSxk72oms354MFwkcSalgeiRR
wnLPC7A2esT/qphfXMFJdPkaTPccZM7rXxkK4nBFb9jz2mTjwyaxUMM23ivrWZzNCfa6wixZ301A
6/RZW5sw6kkY2iToaqzlU/ECraTESxtm/JGxSE+EsTavOSD6FRnc6FZOuW+RrZPz2nBEc96VFtAu
rRMlvz64cdZTZcjK3UyuwwTaVLOgcILmt/v0H/2EFcIYo8hQOU/gFnaJb5xlkPno6OV3MtRLf6vq
vTw2DRGXWmeeLRlX2w5G945rr0w689TWdsjKzODdnoLz4TcPXNYTSCCRRynI7kR3Yodn7mm/XIXI
fPsKg4i1xbGA/If0HkjdMG5xEoCgb9zQFcPILAi/eP28u88KrK18wCDcTTECN6zKr8oiyuQLJ8gg
0/O3nLE8GRleJzBQSaNfgGu9E02P+JLoPfmYpU1tvD9mM2+cVcxhWHw+ggsaYoBAICLeVeur5bKV
v+H1OxdfgWY2WpW2v5m3u8NZ6kiiGsWvKcRqDJUQWrCnWBcNRAtZoykoeKxJU8Xn51g4QRJLW7lW
EE0zVBi9hn7+cKycQoEXvkHr3bM82rj+OHsZnM8iGeEC5u28BGl/cCJ/QNf3lsLDKW9OzY/d9R9C
+aul8j86tv2ITiiZDINLGj4wZeCQrY9JBePH6c1p+R+Fiu097CHG0MejrKCXd755Rb7fBCNn0tRf
li3UvmKhhpIwnHjqK7lRFBKujcprTBBgZ5vcdWbrYZsz4fs9g+xfQkMcbtrtdkadheq2FvqX0X5p
CRI4Fi2iZDQhSwTFQsxfL4dKgNBhoRErtpxpaNMCj8lYeQ7qom6dp7SlkxFxW9kFvIRztR7gcMnu
Vo9/npnaNiPWjhN0OrYvjTADenxmAXI59gnqFbnqyLz/0cod4usxvKiN8c2DikwcQo2Oeutlg9v2
GQOrWvPwsfqpDeqO13izB9O+tqBvQWXQXbkl3lKecV2dSny1N+TnlMibrhdUvlZyv7du8OQ5tyir
1rA7uyxklnuL+XJwoC1ye95wX4JoMxcyTSbYw6PkoyYpbWPT+fcwX4o4emULH2GSYzoCPva3/pbt
GzyB+P7VGqbmW46jyvpUi7/tImh/I9DDsP2aU6osuxzbEO/Sjipk3XuPdg3C4Iq1E1g3+9gj64G0
948+yBALWLi1l2b5bJTO5Tkqp3qGc0BHGQil0yJiv6IP0SobbK1Kk7EktwX8twJDwS3/2MR6LURa
OBMfeIgefcv/cr1B4aUZOW5MO0+jBCXb4htpyl313VXeNFHjpBT2ovCi7APca1OJjrXjbXRYayno
cJtom1F2+tEcdLdcQSaMfbUx53UAPvV8oxalq4pna2Lo1ja/gVTNMULuDqN9i+13jgYD/QNZi9xR
JRQN2m7zSL5lDWhCIXPmP8mQ0hweNxlpykAkMuDX5SCT8uds3fO8LKc2C8kfl8HJ0Ewiz4BH2PVP
zGmKMWLCOCg4NSx0KjEI17XHz631taRoagZA6IGML87EOPlDosKEMtqiMjdvNsR641Z11tGHJurF
a0VoOtFtbCd4rtFlT5TSPnptrGt85vhUs1QiMr+YlBK5u0IrAzRs99hezx1ypTted2CPbTC7Kx7s
h+hTuEzLIeXsjD6xQOkHRDLMgfv+goWZWXU5PSwWwXIOIYQ1s//XmPfY0gt1K9ui7WohjvqUHzPQ
PhYLB930B9zIiGa02m2QxOdzpCvWV6n8MTHCbmN/9aPBMtqB6HK2XILuOpkPoRib7dyxyAzd1R/m
yx1LKxzQZIMUnDvrA9do4x29HyDoSjVs6JLClTaZ2EyOVJ0RTiuxErHjDd5a3r2ltw9VNrtJLlxq
QBOmyUhrJzcv0sQ0DoXAhGBGivZSBKlnIjExKaMqpZa/jtg7v2SO0LO1xJ63t64aZCafrWkpXRC2
5+AbCuoisidcLGoGgoIhqRjbEWobFyAa1XEuRjGOWKnTtZGm6WLD9arj5LeK/PhubxRybSVUlnCK
RFPR+sBMgVJ8INyK5bhzv9EAiiXvosPC01Ls920RSBVLDcuG/AQXBU15EEZhs1rMLNy5l3sAhYcn
qNuY99vfPZNRrGCpDD7TNW5VkTT3ip49E81NVGPa2i6kCRSRz8CP08CgrDglnmiOXNL0Pg6c5bHT
Yp3eg8UF+B3haZREZCB85WB63EiPpTmxkUXuaX+/zHNJucH1PQHl0XqoiT5yoLniJ1HFrvObhCI7
jfeRrS3PBwXKoexcSmEb13PbjJlzGdhTrEEknzYNZEgnFLpbSpp+i21vV4P0yLYHXjqCVIVQa6Xs
FZ42Ns7cg9XDY3dWSySuHWAnckvs8NlP/kAInAbMmKXIsZQfHFdyFngVWInffDdqTOs1pTMKE+Us
5eRCjc9O63QWssT0Ri/5zxWf5oTkWj8z9wZ6kww+UcREQRhHJKcYjkfCO11fKLQ8C0RYGLP5LOGT
jRWEBpHTtLCNW045XYkOghiCzUA8TGp7qFqTFys9RnRCcHqYmtHOZVYqLpdTihpdiQWJmQBUMqLw
Mnnip3i+9UEAOfiMylVNBug63F1TRRezXPyM2o70+vCuN9eJn1PkkuXwPbG2G9o9vt0f0FB5XaLu
QuCNcN84OTTNbvsulAfnc/RrluBwknT56A9JQvQG3CYcuqBC2lNCrh4vBSZfeIXa7ZGcExuA+W3G
PBYnf2s4iAPze0whWCf/+Ee73OfVdMRNM6SUPceUjK+UKADFaf4Qp1b/cOR9/MwV3TMa7iEt242b
KRctco9wiJOSLrYSsS0ruQoZ/BZw3u2/BjKPPOE22jbD6zCbB7wgM0krzGRd4qCY2FNs9/w9Eyia
thP3T+QzVn1DwdmCGu/tNZQavBWrwAi9Lf/jA+GPdnml0qZnOHfwRg+hfHr8Zraby5tTu9V0rmNI
ru0MsxhCHwCbc5o5t+vlpBlqokdAkL+eMy6hh5efFKkr+a1V1K5RzO3BaqXJg0Ph7RAgbmJnMU7H
C8rpzoYT2VH06gX9dOTHGR4UwgdMQ+7dlHe6VFR3dajbIpaMrvG55G2mx3hJoSEDvRmKz36klexR
7Ka7nzxUTsJhePdHKdYOGAw3fp0jT3fITXZGOTwhOuvxe8zgMnEHos82Zr4vCGxUBSpmC/wtL0FJ
xImeO85sMQpsoHCLuMpBa3h/kOC639vPZMMn3Y7qUO9Gw5QAaxQtNy4No/92p89Jlbj898MLsKVV
QojYyqx+OLA/ykSS21whlvwnE+5Yf/zv3ppCktWQWH2ytNEkgFwQHSHnQbjI9aYqCnzoRAT+FfAD
VceFq0LAo9jOuZCCfi42kDOVHgCWf5zoR6AqeBFgWqcYJBdUXDQYroN/wi04OL1Cdomgrio/61mI
C1mIs1DFiLPqWnjYG6kkhcAAzxR3bAHjSpykC+H9MZ/kT8JlZ5fwYWH4fHaU1p7qR6vgd+sHvuCI
20Xc7PWs2zaGN1yZfaBViTUA4/KzctdEQ7uIlp+8OhiDw+xoU2eInt2r5cp8Awk9s/IHZ8PrammF
67y/svos8YFN3QvjQVpeTUzw4T6drNr+3u6NmdYjLbWlhubi+SfAgOPhMbTG4QLlaqOXQU4ysU+l
hoDkk5eAWjFXX4id3+K0HeALIo41sLaIYqjoLla/2LU1rc/HMcGf5FZoNv80CA93H37t9RAJ9K4a
CcE4moIKeNLYJJuc5TdiBWoT3ethSLcyV9+rtkejETFwlaw6GnmNKVr+0BHXm75NAa5N2eUvXFtv
Aum/Ukt3U7n3hhdiIPiPq2Y+YTe0ERMvfeXzqY2k7KqZM4zMy0NP7HkupFHGeGxHxievLFz1axd9
lvppAM+9G5EyleuQJUD0LEVdaad5sQaPY19JP4pOjGU4V4GCYpgcuIVZFmP03xHnG+NCtXkPEjEi
YFt2VzY4gzIOFgIxRtgTVlLsFN3CZ7xUKHrPtXmW0qRlbFCLwQAO1Bt8AbNGuCA/Vw7bDZ6eUXQq
fAW+G+ivStDg2YbttLb5run5Z9DGzEpmgaize/30YaMfCu9z3UrjYUk+spgbse29mw2RuhhBtTsY
MW3rOBRRMggTn+n84Q2LBt4NSxGb/OKrwqZWEoGOzYEK5BGL3IH/FWSreXAnpgbR453O8c8m/Ht3
KbL0NmGU+FNNvNLkiK2kV3/BdA5iYshjXIAS6IAj3t2hxa0xE9rakCewkwFCOHF7W0wiKBKdZ9kV
DmDEdYL9mErou9eahUv+ArC19QhRIKE6glxWsvXv6iJKrglXAF5+PmmIJWK1+ay17A7J/U9aKjZo
Eo543FitMUY6iFAhvWhXse1qPn0P/KmUfL3l67vwYCnn+wMjkrRq4zvT8g4MtQX0WBSBZcPYNVcW
wtK8iMx4JYU/EZsZ2w/oFFZsQ3kicKAe9yhdg/tJHgn7yxepBHYKAhvprzgZ7MDVPHfVQPXtP0ca
EaYNYWcleMTwtSHYPmha4R5ppfRpfqwUVZDNQzPd/sDj6WlTb4pwfFkfdHi9DJOyqKRFwUWRk3nQ
weAWb1BtdeyTuMItunA1pZB1xi5cvpgISoaBSojdMVEgkUGsVvD5MBza9yq5R1g+CEJpkWb+ozPK
YV82nCDsX7jqEO7tRqtRSBqRqAVPUm8n/5QWMuUwZSu6tITc78Z6q0My39Qz3eTeX7/n1T3WD1hX
hXc7ZC1TzvvWytR8O/rmPsIZ1iphPA7IIVi0WmOjxdnns5tduBN+pv3xVN2+N1D9w/nhWc9iAxGr
70dkoZLNQtL1vCzNqthhZBcUQX8FHWcypBJYwFvAhyHCzphHCjN+DwK4QFvWeFHiLkxp42c1r1V9
xyydqH2VccVbSC03V8h1+vLykhXrKjkeKWQZzyYERBl/kaI16/jE9qxt3WiTwey6ySxMZLA2G/lm
UgWeW/Emg18aRYrOKp3Cy7VJlMeNqfsQY87OVlX+2itAVtIAP1KbZZDwWbBEGaX8UDAWpjXceM32
ShNLWiaZQ3HQjMeWySByQxjNNbKAWF75IngKUN8RfUqtajNmMoo3maa0L5+0MkCQzOMknW6c1zwO
F7uDLptL7CiwLfJCEYqn32INxYDhxLmFf6FM2M0rMzMQqW5dtCdM9e8Voxi2Bx0LUIPsqj1ovjrL
CXJiN+S6F3dNxBGcezUKFLkX8bLKRi8yN98v1/eSztLPv9B5zd58tXjpQb+qeum2tTxD+CFkJUw1
QyfBa6Lo3KMZtww/TgKn0d5zPHvtjjtWuR8w1KCQpo2B/4M1zBvTh/HEaVgm7DUeQ6Hg9JMNidf+
XixAUxPT51A1/dUr1Yh+O6qZqaT+dGxNglWIZ4UI38z9Fkm6XP48TGKmuzm8dYRUppF50VvMPjMq
mtF69zvdgap4KGiwf4vOssAs1lGkrLpbm6A8sepS2waO6vP69RqkBUH3mkE4AmanpB8jdrOsEvg+
X+Xfvo+CqdB8forFv/tXxiZm4QgoACJgIUjtmG0hMzmeNbDIMPjjkMeP2AxCWA0jsw2ytDOuOynG
siLbgA8oLKjZeGFxuy/OxKwJr5SFxkqSav/cANCSIeVK1TN8LLCrkHVJHZq4umCMaFt/YCc9X/kB
MI8ugJBao6Ho5DEUNKBOXPBeZLPSdohKjH3e32Tjz4ieYiUDYv0B+9rBNgCEtD7YkdKLo4v8WyqH
tPjjF0hUUzbNGhe2yuG6zRBsvjYLHqHTiGyO2GrW4CsqAlzGov9WPYubQdjSlY1grT2BMnkwZQpS
gIiREVgM1CfphEPD7X6FeCuHApL0HZh1i9+7K5urUNrB5+1kKaeucgC63Q6IhCRfsMAnjb4f45Fe
QIshI+EKNVu/M1kirX6EL23GONCNRpGi/JFCQpP3EYbPmDrOSkxcyUBYgf7Pwhj0PawdM8cNo/On
FPRFiRXLtr9F/1uhOO7ezynM6Ou9ISVWMe11FxiGB+QknQ0U0EDTFh+ltGZPTnK8cCgb5pnkrlJ2
pESDO2lwKbJgZz+E6sN45Vn6XzOu1RdNSlguFLped+XS+Lzb4OI5IBh+CXaD365bNfjXYTfWSev7
N4YC43GJxSO92Ps/PXd3RK20Yud9UCs0C6qPo9PdDI86bBuzw6yHOIgtt1wBWl/H2YyEqxs27JSN
DUcAdh+6eAfExpUyP8MI3FuOSBirDePJKK4MrWG68Xcdq9+V1zibE6maTLMuSe6lR3Q657Ji24iv
AcCpIBGnhSFyr1SlfTZNn9UUf23qOK/g258EVkuDGLsOWZ2Jpi4vDt/D/DsS88EBdubI0bwegx26
GosnZvj+9wbNBTTJKpGcXg4KJqNer+ITaPZFHmbTp7P/U/NKJ1vRfBPzdTM5/XPbZGT/kZ/5Bv8i
fzMD9cQndCaOGEyeqwlNYGJDnSrqfV/PpOONIn9fnDPvyizmeVg7APAe1rpmFncBKxTQ+ZS+khAi
oIIW17btOjNQgtmKTgA2sTITs9cz7eg8lqDnBD4zsTMFZUrvhqLSlZMocTa1ZYK42xzEmvZ1lmGD
ILwyJBGXM2ANKMmMu5FJzCPTrO9+aQrcorOT9QZ10kCsMP3Ln/WBYXrnIQbIdcix+uFzY0qQw+th
n2tmuwCXPkAkhNCuAtxWSUM4bZzEgqBmxettpe5v9ganDb+CxqNI9KPfAHEqa37H2MVieMnBB5FG
nABQDVYtUjbgAJ5godu8jbuqpkfgjHr7f5iYhJpY9qVGPrxWHFdwe7Dj9q2X9BHYplOPA4Ntt6UW
7kEBV8JH2l7hHdKB6ObMWwiAjSasH7RrqQlyrQRR5mMOrkbeGUeqYNrH6hNxKm8zuK98cf6g+Ijy
JtUtqHCnuU7h0GdevRdRso9/NFiVAuWcAo3VKml/1KdknWnrlJqbu5STgsplaVyIh4+pGWvmLbk0
V4JG8mXXvzn//RSbiw56VICsZku0XcH1vinG+skVvgTS2SIbzC6YLr0ZsjZ7Rf1YJ/VP9RyPEvyw
Hj4sLPmKr+dYSRvHXGBLaPR1ncRUMZz/1Q8Uhd5etFx9pv/E4omgbMuC29Vp4xdZkIAlsf+ve346
oZHmbkkc6Ez9B6UL+dzsi9KG0zjDe9NM6fIJ5dn39xyAZRI8bjn5ZujExvECLGZ1DvhB1tiL32rO
ZH7zC3SBzLILSoh6qMFFKX/UdJ7wpBlubldsxktKya6gTjFKU7NDMi4yTLNbKiI5xH0kPcIn8QdP
v9kHzPdsPyrvOpS2vjE2WvFcvEmSjXRVcYoErgvFu7WtQLPtqaqS4zJ8aXAokISNCDpbd0Wmlt86
GK7WTd6zlPil5qRu9VxeUK7zuVk6lVs1ZSHroEqPEbuT7mWlc0v2yoqpdDGETUj4Y2PncNky2qbI
SXjWwd2tcy9EkJW6Uv2LAaNWf8Otb2ba4LgvqEKC6H5RTY0QgWrbH1jGO8bIa8dbTRPlJP79LzTs
7ggUlWfIgN/QBbJBC6TJlR8t1seMxzluAlMeWLe87BRZ8Y67pcQ4on8vlRlrDJPGzrfSScwAZnFg
s5LXlC0SLSyR3gR2/lrK/7EZlAmkGUuHn7VaEVfanQZIypbvZan3Wu5PjvB5EjwEwFL69MaiF6EO
Y34M1i8M0JUZMKN9KZaBFXbUjS2GkIIa/hfPtz+7Q2hRQL1A5DZ23q9X8nbAsC+kndnnbwk7D2J8
VCtP7fIuNnq9z8RF59mhq8SNXES98Q5uuSuFMh2z2jN91rbBEmB73ylEHCBw6+N5OAqVFk2bVTeJ
mswx+4gMUukBw+KGuMbGB6bOhIvoj5gexkj2AiBXxoqSBrn/EUPWlje3DBKHSNdaQf5oqZWUsBRB
uC9uqI2rHaecKGF1eG/+qX7mVfMpgPoesLk8hWlEG0uKynX3JGjdyY0rGHN1uYZ3qREX33Hrf99L
CmHo3xDxPtYl6qKpIoXETF4VzYl1mOkRaqxfdgV/+scExPL6CU0mCBVkZoF/ZW/ZHGbQFDU3QBXw
+nPUNeb1wgHziswpBZAlAyl0cb9RFWaTJxviKr6N1WudvDxeV0B5h6iPc2YskA0OEBXcZRXxT1pf
QzJe/lBgra82KaVIveaCVNPaHQ5/UxjYPhyWXLmnCd4g14P7jU97mQAd37FJXP1IcUoQE5oJOtnN
m5l3kFtgEpGSUBJ+m9yr5LrBpIqu60wvPaUVkLcaypRz+TA4XKa+hodgtmJjE3avBY1tsjXmuDS6
3q6UeZABl4A/1sAhHVX4hqCnn4nGcqnPPNUnNTBjGfuhIPvZ4/KbdDEBHBWRIW700xCgeJVE0iL6
RY2nx/ZXXXUYtneCAMpcEFm+xHerKRAUBFFIoG0CvR57W1/E38XDWLl0KADTXrTI6fomybcQ6hyV
aZu4PeiPE4wqH40/5nt05BtaCSU4hhhD3PAJ7/HhSbgjp9UJfoj7OhI/UuYjiAsDZ73a/E8rrE65
wh6p/xSspUr4r7Nm0but1Vng70Fu/uASf5YuYMM860fczn/s4GcJe1eqRJYRRS3r5avDy9YHcqY9
05hCI7Tj2dW5ibXXsQYTQzZCLt7JafG52K4buMIeju2D9fRazRK3j/5CfEBqQ7HWn8obJsBBRo2W
FOI0F+vn93+FV9aduJ+jjKoxthLiov81F+3IkZjM1GSxnaejDEKCukSes9ST7FeTNaEBVIvBpMDW
fp6EwbuyIR2YRB6qYfj1FYORgq+YJAeYP6sxzEHYjWmOQTzHCByYq90frb8x/ZY79XH79KFJPI1B
IDCy2FKEvOhyMCwMcMntwrL9CEcYG1eBrxOgPl5C0wXnIgg1r0HvXDPKWDpYmNfEH5WWIwDTU8iM
QGPkERy606pvz8LSeRcsDSeMGz3kIQfHt+XEhcCAYZiSYyxtwJY6gCGadwW2cj5gioXkrvNr89Oh
pllmG7XmblXhz+p7MxzJ6Ejre9IVQXFSZtQN6/7C3fP3ftMHVPsPIwsNPW91tlZc/XdiQehK7wVw
Evs0E1It39wkMhJUllQM5v3mprvfVIdBD9GkCQ171Ctp7FNJgf7WElN3hsRzOW7B9gtUoFb3SmI1
zkthtueCB0JFpdh3JBraLcBrekQ/3fqRbyFLY5QC3f6nSNCg/n7+uKWS0sGYaoJYaPU8BmJjClLb
9rK1Kg32uYyJltu92s2VGIrlS45tuG/h0A4GFg77mFLduR+tjToHCtVTmOBGNRY28nejNo4Jha1S
LAWmoubLblXUOag2x/DlF+7h3J+s1uDwE0rHwD6fMHy5QsMMrOwHz3iKgSt7iUu44beK9Vs0s7ow
RaG82jzEuzTL/h+5w23Kx4vab9wFPcSCi7L2OmC33ee9qBa67I/JxroiO9aVImDwvMaYzb8laFqQ
ZrnW88DrJ8+wB1GFVzZLOdJgOAV+vAXw1Dkv05e6BM7HsZuycJOJgsYazDBVuO/Qj8khAYtvWn42
3sCDKqnd0v6IeaSrTLKHY2waedxAkh732C8bTN7qbtpzxFT014oE/Q38qbxHk88rAxl/WLHMQkWg
69jJnuDsLm5+5YfLO4r0yMdm86cOi9X202oUYOxr3haKDikJIvMwK4t5zgvzfz8/SckxPQctsMu6
lQ1doZTfVsqtF8K1xIqKUCQjGyy7kqEN2YCMD7AZaixuIwRGd+GSsqyPD/n2RCIoR/UBRX7DJJgJ
bYMSAEAJJ62x0ENZ5jeBpfWAFOHDJGii5tG2X0ynJtwVzuiiCEfvdkxdOoDII5vLRQzC4nYOMaA0
WfVgHMKz90OLrDBBr0/gRw5aavrJP7fpIxXe0NrakN3W+qzO4Idnzvz007cnUm42yELxcy8cZp2L
if1LCLVrUlmcq58VjDKN3oe2itNCRW0UmTYj+/ZhZt6ZM7IVgVy5T40mDBNR7e1drz9YPkcULieg
wDpLOuV5mgz79VmhK3eEzqGBWu4ycataZT+bz6irA/POyNzX4yVZdnrn05lhjpxFFRTEJm9IfLkV
Mmz3NMOFRl8eAlTrMIEmWgRDuJTTOf/E1AN8hkZ17R22rISlE0GyyW7lXnWg/M9ntENqq3x1mEjj
s513tLxhxRTCp4nfSJyTI153xEXtaZKWrO0w/xYt2HP+++9WU5iIc/Doa0UFa4iy3Ig4Gv/n2/Jj
qhvRiawDxpjiqJcWfuL1qB/Uoh3csGMZ6mnR8MN1OKqtQ2SRm/lccyUKqk+PvE0e6y4JyTd3Z64W
CiMVravseXbbcZ4w4kg+mcw9AQHCIp4k0Z3LFIfSvIAaKc340i9cRYFwpkQ57PTxhpe7HYX2JXWZ
W0NuPfVDnKtzEitMOIeCSE3Yih2M75N5PCUwXvwAtoeDCNa9bcAS7FclKgexk98ONhwE84Vv5OBn
gp58LlTMpvNwfBd62y4vBXQfBmhKTjw/J4RFKUdTCPY1a9NdY1ShGwGBKlfujBaj4A93E9rFnVSR
hQ+XkYVldlNLlfnL2MUKzHlsLNuQYxtLyosOaGVXAU7qAPkSHrx93yEl4OWc7RUjgsEJPYCjZvTj
I6Aet2S+QZC64yBgmXz6tuHzy1FtxnSeRuCSkKfn+/thJdjMQWMWWI6J2vvCfkhfjblVGquBTvsq
2G2jWYa1ju8ds1EWToMaDFb0wEXgltrwCrwKMkD98KkFvmFxbLI42yQzz0pacNX6aS4rU7BFKs7g
6A0EFiFFGJp3coE7Ud0tjxDoTqImubrVa4gmlM3Guxobf0L9SH5BX1vjWl0+WJzTA12sA1quH8UF
zv4nL6yqv4PE/1FTT5a+Euefwi23Vt/5Y5t7a8ZPhYdHISj/j48BYsRTmQnFsz4F+sm92T2GBYuB
Qk00c63BvL22EWKaXP3+iBEOh58RhrtrKyKDeTa1Gp1iRP67SLrbU42l60UZDfYBHDQYD8SqTmx9
C2EC7OJpWSpZIeOT14eCy7ED/MC4RCFqLoKi3sgHQuRt01JiHPIZ21cS/zljmLEpoAVLvfTS3hPc
Mnfti65lGw9ZkC3mOY/BbAvC1+vSLbmmgUYahfTLaD5JIaEf3wkVzA4pmcATbVWGawAdYfDod5G6
WWbx0pQb4Ii0rqsYPI7OEeDAYiJL+2QQC24sl9XHAHYhEd1KVnlAUHxQ68hDynd5aOIaQL76XMi7
wGaj8VHC/i5Zun0sPHHY4tHAJSzmph9RahRXt17DFt0rvG8bx7MEV/zpcGt3EPfKHumR4IBf4wLA
qz48+9Zlh9XalYdllOAty4mnZn+PfCN77U/lBB+3coSMm57tY4M3v4wnmWSsVeB3CvP49uYKkwTa
M6+RooDA4pfBtXddIfUdh+Zeq1CN66B6hGAuTg6tJANu3Q0GcBngIfKgnHiv+65FH9OQxm5F7ZW5
G9UyuexQ7lfu5UnQC3FARMsPBpePKeww+vWt+8f/5oqxi58on9b9KtnNhHbvI3zcG0EmR5ZdnY6W
d5nqbVMh9EB4DjRdkC+v2HgREXZ6sdRdW9EwRS5FEn9YSaeACeB1HHbuYCiMd8jiI5A/AFCvyMOc
tZyJX+EY9DiGoTLdIAyzJ6tvC+2BoP1XcE+kbuC6/P77Xxbj+FQ/+0h1VgjlOUgWTimuf5EvkpUa
1upvrWgmEJvf9JZdZj1z5FdtkaRRXKFBaMxeKcIIoUs8B2kbGsfPifsb3bt47+Lx+zclVqPCK5AP
WEwlGJP5dCCGmYlaAT3dL5kgL0mAxOSZAke4wen8gDxFrrgIT2w9lEpEQMvf/H3OkBnYa6g/Sla1
qb4d9VAxRG0OXWICsBHhkNGEQZSAWN56VZRQ1t78TF1ykdb2STK6Hl8FApV4jQclQcCwLFvccgvN
+ind9Bxa6W9/MWITFTWaQLYFyB3tNjcG7/Zma/HMyM+EEYkTmAVhY4It6C18X2CvoQyGkQRCEogi
Xab+yT6KR+ON6g6vhO5AjZ/7M0VtnlIzFmhRNv3bMg90aCelEGccgPZOo/cDJgaTysb6Ua329kAl
nJ42vcjWUOL/Tch7OnhMO1TGCfHMs7qBRjeUPU8jivlqHrrX3xDlQhrIQhXa7vQIVy80ReSd/W+9
/LcHQJtQMVoh8a7MPvzvQcfNGym+HP41a3D6OwZYs349M8EaMoPQ8TA005xQhuhlrXkbwu2j6xP1
9G614zeEbk/04CHbph+cAB/LIfjpfc2oYI+nwp/qizDt6ZWJfzXdLiunYcaFZzJRxAYtUjK8cE4P
vhupVmGzU/wMzc8qUyq6VNzBJYn+UJmd0SeyV2rkp0HVQUAplwHfe8xr8YByAYFTJ7LP16Fu3pAr
8NsKa8cx1+Q2lw7ZVbNLs8z4ibI6so9YZmFVPuE9SdQkyfXlo77AAQfXCjGjHvC9Mi6weutb+2yQ
JogBdxl2EOxykbF+5TjwmuM7QyC4qA2s/cGj5cY4iLPaXDTlO5VeIYMWNhOCizfWrfvu1nWMP0TA
uQ4S6ZQIz7fgjNy99Codm0kgkJtqdLUXW2VlwcpT4ioBKE9BlXKjgSKEXL9Ee26sqUN/BfYmN+6V
fr0bF/TgTMJ0fsViE2qASl1ir+KPai2zj1Op6KTnDhNq9lvxjVD6SxnTDhVjLWmvi5wkD32dRkLJ
BAvQK6y9ON0PZgKoUj2HS/+vT//2bDqH+ZrUN8VPFCZl9prClcVM8cAyQN/y1kLRHTTTMs5+eZPB
aQEHh5zLJf86Pee07tfDwFoPUjToCxIcBs5/Eyaq5d0YWdp1j8T2nhcH2Gf36NBhzY3kfDldj5F6
FIE4m1OKrxfH/duqgIohujgw33r0fv8A+5NFQ47EGGI7vcDOUoLS3BP8+qZ8DTONQL2PDNdKxqQc
CNfAfXdOE/GZP+OI9bsd2bJBzF3Z6ieZKoCVXvapyxasDWUIMi99l2Z5pcLcNMu5ns2TPN13pdu4
IG58Ft1RMjdCzncHq3XZwWezkzeCzAJYA+xU37eOVxNxG9bWuhKdRP/hV13EfYYHHP4a1UDQROn+
8cu+o876O7yM2fIdf43Sf4PLQ/WHCULC+q+XKhh9eDSacvYj4PK88W1FPyrkoMqYqqYNNvAtAyJe
B5HxismlUg7AZneO5DW76m3mJQQlLwcFIYFOIp8N4E/kVdp19+tF9dxFF/k+Xet+8IyHbOUCXECO
jBpLyn3KWgu5b8b2uFci/7LTy+fNVZe0lpRK/hg8WhpCpzOLgIR4AtaH4abMmB4aFbFNdT/NQI9H
tmbVX7Lx54oFo4jTnWMWNy7pp1azwoSP+l6zKiCujDKv10ubQDmvvgFT2SWCWQFjuwvea8doot0k
xXUuB0HtjcDTqDXF3H36QTBaxLfjmHgRgOsPOffs05ZEusgRixJeGHyDRISqCrcnU5PSqYQeHYb+
Wcfxtc6Z0gE4skfK2nLIj9PuzwFY14g43jS8Dx/hIS6nBp5i4iuuCIIKbBOOZXKANw4BnfNavnvX
2uRx9TsNrk12s4L4c5yjKIvrffBVe4Vby9SMZu0MkonqnTabSaF3hypHGJve/PPNv9Iy0FyenF0u
BYzbP1sHlAJROBXsCmuWuSVhI/NvnhxZeBUfXd/7wB35eeZ+NYIBqiqJXCGfEYXaxUYrADbviQYi
kn7oswBRJBiIcz/J8osnf6cuGH2eZlC5/uy+5tL2BkgPOMN42Bjmjo3TtclFfuCqhwLOcyW9TX0w
fCt5p6B01bVEHocfWsgwirksdZlL+NO9PMijMkChplpDE/AY3jKFSJ/3+TsIlzxavkDQ25jrNbVV
GCSx5XpogU/B4/1YleTJ2B9f5ePwwVQ4IkkFwDOu7JdhaSMISQ7anM2uhKArLLW5ev1m+qlnfXqW
n2p9HsCidA3TX8W+x3OU+I8847SQEQKnt6HlG4pX6X2eEvoxAXH2mDb8mMxHKZBHTMrO/Eqa4gP4
xxcXbq/W51duMns498//Xlr74UPmlbhXGUXqfyxn7kGhgd5EEVCWfT0OJeztdJKyvvAYv0Y3orA0
EWxjjxQeDF1mDSqDas1hJKkaOy350/p3m9gpUCguuzO08wPVlR2rF57DUeflULF59NDDZzx3oj7a
ayG2l3AQImUkcqiL+sjY6osZV4nrfJxCxfpzx9ExKqafjRbObLyQS/jZ/pyhK+zu/D2q16D0HP14
9iG58g3pGDrhrr5SlPhu2sTeSfhsuuXJjniiSNzlOg3tyeBwq27NthH2yJgW/PNt6AFtsvK0R2Dv
Gtw6/5FkGrRcxUmo9u4cA7Rs2jBizkANPD5EmBdMjKJ+HwIQXPC0nbSzPw53554eufngrGrNPbo7
dF8IjzY0UxeAc/jE/1QEhjiibMgLkvUjLgDE4/QXTphSaEH5TaZNSHdUsVMUVw+3shJST0CkI7VE
Fo0GyN+KInXn9x70ZIm55j5V5C2STQCvXjLIlAO9LaPUO867YWdALUkwQ3YtkyzqtxVULvq5sqWP
E8qDRF2sN/FSjybXQ4/c9xjmpknX/WFUSU3YL9risS2EfQs3zdZ47hukkLkd9G6IJZDIdH1ngzRg
8n5x6qdmDIMlHYymKs2fVxzxHy2wzSazg1eiJbp98MYGJiBLRoATLliUCseQiVWPzFuicdjMuPMx
yTlKy5l3PRFCwOzV1yrEYDDAlb+FwmLbbMhZibcX1tu0lLputmq5Hypow43zNJqtsk/N28+H2LTW
Qx3tLKtTvma+HM18ql7chGBIIjTCGCM9aYpuiWdlIBYa/Z5Kw2PdFg3jYMhZ5sz+uL6kI53klyHW
ZQcmL43W8y66pWvD3X/+hDeJVHXiD2iWK+c+XMzE4cOJPW8c+pgv32l0UIZOEJ0vAmMOsE3r/0eT
xrTkJcC8LiEer5HH66ZWOnHyCPidNErNx2gtg1hXJZEKS0z5y1Nl96hFTispLvhiR91FwfDd2nb0
0/Q3i3xdPCmb1HIjfzYjmbUScL6RUFlN05Mb2jpASoxeCF7hdFjmd/5mcE2k48Sh+SrXeVmRxbMY
ZOna5yEQLjDlIq0avI8Wy8/2kOLDytx82go8ehL0ZyhZMjTFP6qLj0uf5cDXV43kQ9jTBiI0RSV9
vAGciUDr8SIx+fqK8Qg9pL9V9HtLjO4O9UuLfDNH1eQk6AjnWC4aMBM2YpfFeiUIs6lP9xQvGeSf
MYr1jyzYzV7KNzNCpWOmmTdBPDElCsfbnVKEzYNCdcCsaCSHJYwc5TGrI7VYavF8e+vaYi1YwwUQ
1I0lXyzRFo74cIkIFYpH7l1+6P1nNDDhZGLAiYQRe//s2UhxgnDx+AkfYMhXGMsRXomudlvL99IU
7I/HMz/cfJ1RPa6v2nLkL6DVtRqWeSdfydZ7d+NOuxE0d4exaCNyhpbw6oA2b5mx7OrdK/PVFaXZ
GDxjJqDF5sCBbJPVMn8uVxq779Zf6rGtRs0FxCKoz0uXmkveUcIsutJ7M40ZxlXyS4tJRlhAVF+E
lzmBWUa3bLVWxJKfunmdHPu2b2hyzYwZsk5j7h031TWH56AqjGoHyRGVsVHMDbHyKhYjyLJE7jOx
Es+dz1wLz8PRHayJ1LTOSFx1yGS4REVOkymz/4gv07t6hWlN6BzRvFVRtvMbkcKX4BvPq0OqcoO4
B2HJ6Gl1BOdGBG78Sn5AUscevf+B+m8ua29lo8rgZmm3RyOTSdJhJBVzIwox6JDRwP8A7MFnz0aJ
imMVoGyp8NI3bmESF3aJxSkySJA9TWXDp612WwTgDq/9x/HnvpNUL68AGCHtfydWbXWg8jBBHGBz
VAjDr0v9DQOyRmXdF7DmiLjlm7FambpEnsozjii6njcU2vpRqmx2TMl+lhbBHssUbtkwQGNIscCI
US34xyCcWLyGvsEbVG8In87ILPqExj7uYaHCGpAPJdQbiartlTEfSKU9piMY/cQzUcpjcYYG7+yx
Veed/Ptr1cGYkk+c5c6XS6IAxRj03H+e3TUtjuauOLqtgup9RRHLiOpgUY9gg2412lOBPl5jS0Rn
1Q2F65J1bPHfATZhs/fZLesgpr5rWaIFOFwVVologIyK0QQH0xMeIu98lIzEaeL72yZq7sNJ/THo
8HdCnpXtF8hECLEGNk7TiwwktSdkqhTeVIveEYNmAUOuKWkq75cet9VT61nvzMA3P860hbcvGKkO
sbcz/ULdVdAFXEUWCfquVsv5X9yEFWR3YGig2yIDT/KAlNoGy2U41MOvzUi/6aRJf/wYAIa/Ibdg
9hTD0FslX7A9uP9+Q8LRMKDcBgpw87N6MWLBlBGUSxSMd5kXg5eceSVVXl/ttX214197VxCbXZ/C
MqfxRdhOitAOtuZk+5u8PRD/USH/Fx/Az/u9XHX2Go0owYP9TqxPSIyxdyPT8740NOklyQLWBHBM
pfE1DBPq2yEeTouUGqEWioB9Ad6P6W73IWJqKj8jEYlaAWEUGIl9JJfz642wHn5Miv0GwNUvqF9Y
Ss4mh8l4B+dzHKIBeLLpbh2ero7ahDQgRVneHaOhvzBh/2pIqBpaGRnV8BmUTZimS76rZKYsVCBJ
6e2sBANoLpn0vifxe+OvjYBbz/59SPhkW8U8mocWy9cVx66C319D+6whxN/tR6bHHpRefqG3Wziu
epDT8ltW2uHDHQdYRxX/iRHDV2bRu683JjxSHf/uHu13CBNBQkMeH2w+IVZbnMVVK49ftfudLUf6
q4WbNULYyKsMVx9qoovmGxG9ctVgDpkxiQBVm/RE4UYYtlH3F0b/iohkLpohpEPRLyKgvh2acTM1
LK6z1QfS/XxjxTGY8zPszPceVq+YRU2p2vCqBoJPOplSstYXIk4FYUoy//w6gTiC33iZ0z5jtl1A
y7kThXCKk4MbzWK+QTCo9Go5O4RCFj7WNt1RF9GXlL0+rjU42PXojLkezKkInKqmQOCA1bqY13bM
PvyhX4foYoHEpPULncelwj6VgS6Y0tQEcPpYP4QmObF+DvglLtKCi3XG70CVOQPwrGR/iy887PJd
bh9nMhn/CVEjoVBwvkKYFDd6Jmau2nUII60m2wmFee6FCJ3808GoAKI02pjWIO6Ax+QR2klMmN2U
kaEpIl6vCmHHFRSMIBb5pfTX+Y2vtxYkOxkw1UV5w4re35dLap6aTwJdNaZVVECpYmuVMLFWqIjQ
HXZbT/SZad9Ae2Xsqi0lnsAOb9VlTSaEYHL3Y8P7zgLb9GIsqAuyaofuJtCbPzUnmX6bhxj8MhYS
DAy/j+HDvgL51wK1amntlkAIEp9beciFGxV4zGdD83lRlZBIz89zsfNdUdk9SCn7p0ui9g4XBoTC
/A5QD6qRGfs3wN0Ji4mYah3KHHaz51SiNfr5VBMmTKFlL+693TPBwGS/gwyFA+XUx22gMqdrHS8b
csWw2OxGj3ufWZmMohyFh1xTk+hqGqeyGigt3CgapUEa/owRuW5ha4xKdo9aSs1cNaslVXGP4hAi
JjGcHwljQzCJOwl2iCpxdiQbMmrAIE4DanTPa84xwgfvogAMq6mcFpAfBLYowLkkU1cu+2BLDFUo
oQUorjBkb2uLkwIIKprNC3z7U9lUVH2SsbSgKWq0ZPMD8Llqh1/ezg3MfKkcJl2KlgXaFpGI1YAC
ZyX/Qft743eES7xj0mCrY1PtcKUFeX9MBDeuxgYQZ3JJ+fT4MEvwbyYZOyWfYVPqieTnnGYzrQD4
aFNS1JoobhNVIf6X66yUS3Iw83+/Pxup9PrUo2gieXp1zyjugKNcv5F/7aMGpUpYOuGIQIv+WUFc
aBvQFDPgiPLIDo8+5nh/P30mzDHCZMlcOYb14eIsVTOa9h3K5OvS3PSILI+LxAv51yr+Iu5JaZRj
lXtr5Uz1W4j2BcFyyNEbO/QxU+WMil5Hg+TEihFNvLY8vl5taGbe69ZAkqUOWo1adSPu2Y0TsEIw
SKzWk8klCSZbknBav0Lg8hnGqCo0pDdJVRf2WSEgXIS8JrzofIVe6P5Tm5W2VSq0CjRB01yQBP3i
Y0mrJ8NVdHRlZYK6oawx329UePH0GtYC7fAqAyib4MPt1LDQMmwA3uhkmOkD42nM3fxvshuH8gFm
lrG76YqBRxqnBsGADZI4tO+I5JUgjH0OmOU7K8hWPz0nTAG+RgjlHQO+auaO8rmwNolk6/YH7JM1
OyPISbnVWXIQyVSBiBE6Ubd1Hrvm2Jt+HEjKjKYVbN9sYbE19P8a5cppWu6fcxpQbvRmbHZEcbC5
tFFjQCEw/8/dYnFGriXLckFX3WJMRhFqCMnHxiv7PVuvKLELH+6Stj1kbuoAtwVFYn5aIbH/FY5/
SDQqfPUBSSlKCKzyKcY9I+nwaw2A0wpLzNc3sxvUHHKm+EPpOoSs774keSD9UCGURXL1tIXz7jTe
OTBBck2WG1sIcRQB9rPz54T7Ke9wStNFewd8TLSikdoZ0s7vqEYbJJT9unLRuORNYOvykSOgwKUe
ixbz8eC6mXx7U/cXb/NHaP1CrYWu6XF6u/4IBb9xSP0LD6YjhsA0C4dYLIkirGyvR1fs5GW6GcOe
ybwq+1bncVVOamaVVxQOtUrsEMpBKYZMwMDaKI5p27VfVyQSvzws60NIUwz+KZ5XJvcUPjlgCCEv
wKvFc7iyNKHHi97VcueE8WlUurq/D6IG8EveyhcKBQ8tE+vZo6yN1e5sXK3GrOExelEHpGbWtGG5
elg8YQHVXKKUlTdDTjyFc9/D0/vB4meishARRQH37uopCtM3JhDmkYl7TZEgJv+n2dOfiBnxgrNX
Uth6mxqjhYHGr4ZANKplV7ZYJC3iCGe0HOz8nU58Euy0U+lgqJ8DpnZFcwksFyY3sD79GE/I34k8
yzR93YOZctpiqK1WWkHPE4h8LGIEY4Jg74tALCtlD/KT9orCs9XPw/EZzIYe8vWD82aUotgy7gQv
j1iHZECjCH+SaHCoaefhlF0QMy+F10E9pIu7mSj2MI2gjsLm3qDYEQ58shzcunY2cjuuqUfVbxk6
eYApipDJCN2jqRWQFLF01cckfAsb7br5XASnKGXMXhdiuXkHtoPjyA45yyIIDZ3CkZxKUeYxmrSu
FBx+eYFTGDyEgfG71s9VrybqUJ/4/A82vc2kPYlyNRW8KzLzPu6awOsCiU4ZOmsntU3B+KhX3TDr
vvQwi1BfU+9xpkQT2oBEcLPga/T4XnBMIao7l303mCuZX1NoS0sns9sqbebJq6EUiTfwnciiMbP+
Zi3N99Xw25ttOkbZCMjYDWcNu7a42JIC/C8EL2mwK8soV2M4DK1OwJEjjM9owD3Af2EE23cqiWdw
1/aABAQKLggzqCtPPVs/K7F59Ecyt+RCNUp8XIbgAT+zXMCuOC05QO2km67eoeAnR7vHODGWQMlM
c1BqIUeSqawIqYlarKN2eaRIt713+arwPwQkVbVRM1DRx6SWJqvr+Ha7QefR15lNaVUaYHihQgob
b3a3ZEGIPkLo+j+7oFIwkyCeiauAwDHr1Ojfq1thWSt7xOKfVrmY0UhGR8ETcDUCkA44XtXuivhQ
WfY2r7vQ4BRpNQVUGfVkHA4QE2wUUOdCJ4MzdPMLt7yw9cv5KvMwpxHLpZXfgZ5li9cpvJliMjsg
weD822hWAfBp+c4Se6bQgBPrNurVURUoH4JhtWVdVnQ6JJxpzbMv6uyv5Y3FCtCj/5yZVdIBIekW
lGRB4HmY6k4JCp12QarPN7GgN2MFn15d9prHM11QyRyMSkhfJghsX1wpVNryzQvbBE5rUHAox9IN
E7H8tDAWgt/m0a4NeZqJdzWEkX3ZjGqtJ93hOpWaFGm3tcmRifqwd5LPXeSRrPbUusUh4ZDZcjw3
OiGA4/gcteRRoll6MiUTYIi0ZMwtDvAgrwrPYJGIQDSnQiLnRZ5flMwsmT0/ZYdgphbPPsIpbvn/
DD6IfduOYqF19GyULbiYJJh8hicAVR2aIM7o6YsuQ6uG/XLspq8Svom657J9L8RvhNkWhr/ke8ea
DY6GdwsxqVQIYb3e/GV3qBKNiXkohOibGkCtmFLnO1DGkEeex1i30RjWkpI2ge9s9A7lWYc2PuIQ
03DAOYYDQBZzZ+0qcLmlx4/LrzitcClha7/wvRTQYlKyUZGJ2I9lrj9G7L0zo0FkhOto6kJur3lQ
0s8pEssONobuValmabV30+3nmajc1HVjwTV6ClDntljb2wWqfPRaErsm2C66GXcwFL1smco5krbu
uASrtdyCI5i6Tu236lBQLybSl/vb3QInBwfe5huUQ5hEZNlED7ek80M2y9XVdqFRcRby5NakpV6C
/7LQfyB+fR25B2TlHyH+ni+d4TkBPBomGJDrabMc604I7YqriZASgppm0TTfqGF1WxhZLEQH+oOR
wJmg4LLu3MbTWrvqMse7osqleuxyV+P1L78rR41uuecQMXjHOgb3Mn0cMHVrxHSpvIQSTBV7mFgh
OTPLxEAV8DZ92rB00+SIwlO1Msb4PAIZS5jny4Ku2AxxZw258DEVG1fzGdIPeDJFIITmZdGevLR3
/s+e6GcAx/l3+YW+j50ei2OgzRuGFETe8HtoahVLjc6SiX/KXDLfrQWoJgyfb+5LvFFG9G/NSEpY
lLxxKSP31kyAgU+ayRFjcoJhxGxCHnDDjdw+VXC0qT2i/xkNoOPK/InhGV6zvifsG5QBrhwI4dKd
kL61z6Ivp0xoiHoaun/PzU2IEAf9cADS2xf5hPMH2gwQWrw3swqSSxJnfW8dJn64YiAOkN6gfusQ
FJ2f6w/Rc2089yUIrojjNrhoDLw/+AY7H/klKMo91IS2RtH7/PtnaRMxfZ3o/36em8GZGBYoSSg6
xoD7myX3TgZff99AV4cy7WV3Mn0Y8Kb5FkRqLexBjhyAng0kf8Ie/aCPyY/Djfj7yq0lBmSHWdzY
HQNd1ZqFt/ZhmVcu3YYSwGD4qggKYs8BhHUlXS0K5mcx5nzFDbZAv+7xR01E062r/kMw6CWYjrv7
4YucCwhq2QnFiGZUQINxAJKIuFbAIy3hXG7uOa0mAQFHIycmEEQul1hWf/N23/JqBEaZkqzJ15iW
1B/3eMtDhxZrYbeKSr1hzL9Qnw6VHrZKBrhjvIBTPBfCQ+87RDipCiqTWgtXCTpJ30ZtVs7AQYkF
1/Az7cEmoupWw0udq9yrO5toPJkTl3N5fmvumfJyjUXqp/tW6a61Ne7Sh7VtlSfcxeVfaT1ZRctS
GD+tRRVPqHVeE+YDPTFWCWJ5Sz4n+QjrqmjuwO8M2qZ//HVbrQYJchd1f3Ut6udQIMq+mgw3jGqq
TtBDCkPK6X0r/np66trF3KJZkZ+x0xtxQnApbHSdL+NsalwhPMVM91rPGsM3FjVYAglstce5O7RS
g9EuTm6HQkkYOZPptHZkfaA/cMDlsKZQFJZtkaVSuFoutwLhTa0NrfSckAKUkq1JXKNyPhGPdYZB
L4HGjC3qV7ceOS7n0Sx4IGQ3EMImvCJkP7dPhrjFUhbQmJR0VtmqDCn8enTJtv8hjbIMBUgN9CsC
3lT3AWIxKin3y/v2AxAv7D3HHm+3M1lLBhlD7VEmeEZsfyXO0zROPTZj/YLTJO4YPzB1MD+vPQaE
MacIOnJPiJ9j/1mL+dIEz4EPGTQy90l9NczLgRxhp1vQwUffWqixiojU3tP7eM95HQVR46MxnBOJ
fx/MWxzMWWkIIOYzS5Am6nXLcbHv1DFXWo+nX8j855uaQ/eRepomGzao2rfayZLKxlPYVkhADaSO
10Fr9pVZpolyAszgMekNMTdUkmo+jjSZg/ISrSXOOQt0Mn5HFrvMG6yaqwsH+Ez84FUHD+d2zkIi
yfJsMxALCFqHmEd/Y/vPyU+ACg0fGLVtj4vepHeqPbQ9NxJ2p3qygG8yK1FXDsgyY8Ia/64y2h7B
e16pmJWQ0WiM3qm5SyAFh1H2SbZtsd63tPcDcT+ekhwobQ70xXJl3jogXFhGm4KYFlxTfMV3dW2p
smf/8SkFm0baO0odpOP2vPlkZOkFYiOQuBlF8VF1MrF/3qdO59BAvJtillOmMO71ksR51dkfuacc
TmbgFvHHyHWAB+m3uhLnoDYtW8n3yEBnSfk5WlU/q2EY7iWj5nOXYfxgZeA4iQPaXPvDybar8Qks
WcK3kqdXRm557FYAhh5zcx4EPBUviL80V1IYcRkxQVXl+N87jMlsgnLeJVqg4HuTF11/vPmLDA8p
oMa4FWFX7pTm4/WwaJ7jS22dhGUQtALmJGej+4n+pPuC00NH1jXI8wma2dEtK4CJ2P5GdvWCKxUb
K1qBCwN0NFyuxTztTfIkDYZ22Wysz2ac+3XmymgkGWM6nY17MW8+carF/gbyuo0PwdkxrOTFl22N
xMMpQP8wTDfbFve4OAtWlCaNt5f0VudZw3Z2vJow0byUa3BH8WGGnrfQ1c+RUxdesiN0Y1om4wEj
a5BMTuyjm/B1iJHN/P2neRTt2xYHGT6nF2tiqpXB8kBQkOUxKHdbVrINpWK6LXmQp5XOvVbOXkWA
xU5mcxul//X09Uds05drcZToFUts+kWopG7myCFnjnEJtKkmQ8CliO3Js4q3t0CTKpm8C0+hKkJw
rLfhD9Aa54s5FIb9TulJ3JCF9i2oFO94Qll2nO/BVaPKcBYUSFVBFc5yf7YCKW1lxi6TOUcIitM8
Sesoe+lkyu8Jd29d+WHSj2BJFlP7S8ha7AU/9rqt0t5io9+FM61KEpxyO0lHnFDU10/9BbeRQF6W
f2DVBfSFCINO4kms3uSP1FpWCplkAatwMZs4Gpl7wDols6BzMPZpdlFg4769XQCtSHdYIMh5vij5
XfQBNxM5RjEo38wxjZQROUl454KiEALcvtD8aTUd02uSzQk+VY2iKLPdM67I6k0oAjGWz69nW+kB
iBXx/ArSmC269oIyaWEKCM8EJ4n2OM6xOrD4lQpnQ8XGDGPGNHXIYnhWuBCC/o2G44aeYEbKIqsv
0Ejx5L/PoGJIzOF8pprxsboDacIyNnbchZS10bqHLO4LGUK/hj+OzSn5MqtHq7+lRR6mkPfaLRlZ
cFNEP/QQ2gSvFrJUnoLhELFi4Xsf7B61y76T4g76znrnmHc0REXXE4QTM5tlSKS9JNcxsTJasW2Y
g1PUH3a1t54k3CcP3/RPG4dFWOd0Vy069ppq0Gk4w4NbaNq5mT5tba8TNYP4WuU5tocgUvYtriWo
7Ru7DUhgYDLCHOiW44zM+HVzNsSrPmUtrPigKfOZ7zZqTjEL+dZ19qteuLwfjyd0OC1wOUkTXDlT
TjG8DR8UYJgnDvTi6JTPyGqsYWA3PcHg50wld07QD5km1KK0MxTOnSEWHjHJDUJ3+qG2+yeOrDTQ
N0J6WAjtX0yseE+RNtX9aTGT5+XigykK03PTnwa92lTpGB+vVbzNyYqikOACoiAjKwJ0GwTnIMsf
aFzWA5wKtphkDl/tvYVQPoFWp/1rfa+gW48mHy3qEUYjJ6RxcUxrZqo+RrSVTexTEFUH9CR/ZUin
TLro8FqZFpoCwufA4NTXMKsozSx3N1/Vl1rgSfzSUVx3hhfdkavle5vTaXIZWI/G2jx9zSy6aMLw
IgCRP8iGEJ73YNiyeOWG7qtErnkkRPqba6P0WRhRhpFvWICB9YL+iJPV0Epc2WyCkQGt6YujhPqS
2+p3YIFXNL5dqyzabba+RYa7gO/JwzHyEqypkOX2LRZnh9l0aeta8pDi6gr9m+RqhsCsYTi0cuLw
Lx206fEEFu1/SyceewKk3A8m8paJdlXYWL5w+MG4uNujDgq9sNAa/xQDjMQxvQzsshmqcJpPe+MH
+X3RdmDbNbHqB4Vv9AltEZ1ooNmyNH4/4ROTlrUwxcaABH8ByUw3Oxfj6LS9D6FkwPWmn4trSlmC
yRc9DCjeq3CZJBOmGnIobx8eUK/k0w+gP4VMIMf1oQYeMHO9n/L4zNhbl1pHaBjTkstTMq8Tw+7E
h4PC7GEVGQfXGjwv/fEcmO7BTBwDeyW82aCvVIQYfYa3uR+baiTe3Rh9z6xNfPQ/pT9Et7Bx2DU7
F1fqUeZyMByP5EJbvhiLNfy061yYK9qn4qVKk6Pb17S5hNVEQqw++wg8elKD4mGJojWSsP4LfIMM
2CQdbqkx2lgHTh7ja1bUunvrM3SPRqteJdQ7giz4W5fDR9mvuiPFPzXs3PTqBe1cdvB+iK3TaztN
gYw4caYxY7B/As1Qvf8d0UIsIblWeQxiPUNtRW62uxsM3ThXyjakoCW3FxHuViR8XQhRMOvv6PqN
1eKqkWfj8ckxX66t1MGUGuOtFu2QB4+fU9tly9EsAtlBpsCn1w7xnG4pwJ4Qg1dpvmHSQPj9gpp7
lIjFJwav/5tEnzFsgcaXX9oXzeLSyfzSOqNV4FSYX0VTnzia8/j9Q36Cas1T4IuANCvoF5pHQFqT
eZFWRPy7kH0ugqUCLuLEExvnCBlJ0xAA5hFAMXwS4lOk89U1Ax3w4PhL6PNu3AQPVttIeJI+uQch
99WIbl5WoTT45JEbmF6unOds9J52M2JvQpr11H+e1o3QjaaZ9zwfLBtDMpGcdk8G7OqukJH/+t0h
xVpx3Nxq+CaRakcPDhphK1qhG1zVlmBmEYBdQO8qWlzIghao706fe66JKEGJvnGS/esZh4RC42DY
gs4gAYEuqIHY7QfRA1D5rQ9BnI4E4T3A/iBdyJg9c6XeT5B5NMF+e9ZDhrZmzRFRhIgG11HUxbH5
NCp8vzBGXHKL+RXSQixNieSM00m7sphN7YHNMIIfehliXI+6UXVUHFWPUInGzWCQkpEzyKEnfPhh
JLumEYNBK02OJrEcl7ccSOX/vFbhtxDvgE3ki8cWLUROz4heNo7P1AgHqML/phnHd4QlcgG1FUYZ
iZwf4WEsAKZZIO1yATuTrvjDvSs4pLdv8GB0BE4R0/tdqk8FSFrMaFPv8u9Fw9ttWPEBLZwk11IN
ktGfSfNF5cqSVC4Zf7KGY8/dDbLZC5i8rfNJnoi/KD5HqET+Q231Po39eyOoHfI2MPevT/22dghe
8Bc76fDF8/wg6yWwmWECj07K7bMUj5Wxq8pFkZVKr+jWrhEgVehmsuKcNCgxe9b35ul+1SYPgoWY
oUg7pwrR0SC1DIJ6cc58/oIgXRL4sOftJECUWV27TcncPBSUjQd8Zpvn55vydx49qbPXZ2UZ/PEd
eHBIvn8qyw7o+R4AqvKm91HuofMwWwosbcmZt2qskbjxmCOV0y9XA3l2BHUYyZ058TsV9E1PxM0v
rUtuQI7T77dL23dqytHPgcDGa0g8O5yDKzKQeFi+cRPXjDsSvL1iPyiwepJkPJyLvnTjGMuBpn9W
YaTpPG/4UscSzn6HN6oAgCY1eGE4hXAPlXsOrF7rBnoIBhvkzu/b3PxxT0DZOVLhMEEr3BQg4WQ2
bDAaDt94NNgJtqF2rlm6GGEb9NxOzxaldBtOO8YCS5RoWheF9jMFydF4IzMLnuT7LwJM4JQIjY62
z4GP5Rnmr9lIsHAjmDogVWg9AwPlAnvlCdBWg9JdcwWmIaNVXPvx2X0GqQVarr4Y8JOvh9LGmGL9
w3SW2Oj0QSRnlrKN1/NlSOJBwjmDBjT0+tirEEx/cD6peBekuMSz8y6TsRD2tlWH5hiXOo9XQfrR
zRmQAosYX0mNLfzmxRrTkIggTXRKkhtLMb0vQx7GljyC6znLRnw5kkyEZn7+bhGwxSwh7r70iqiW
KtIgUJkJ8xU+aQtK2D1nq8ZCzobQaFPJ1qtahm0XlPHHmeEzpDCROa5GBC5iCLBuM35AjrQy2Mjk
HAewvviFSJ1Avu9Fj1TO/p9OCyC7AX3YmYurBxWfKW6rxVTNWAw8/mBxoPfKQQG3NfUHuDTbJzEv
d5vDYkBDz6Yd0Ze9G93/U0bwpJSCVyV2T0qi93SUrxAd7V5f0Za6jC7U1f6vk/vE1nm1ttWLXp3d
iM1w3/65BTk/U43Tkp1PmAIxS0cQKL8Fhts0JV7hQOL01xDdOs1HvvYcmkiuqF7SxerDWtuW4rA7
nTWAc2RmZ0W0MtL/W13QStp67NA3ymiUdVoSAzROw/U6+A/D1rWWwZeIltKSvFKILqb6bdfGd5pP
YKXSDfpmF2pDjw3soOuL6cN1tu8rHt+/3M4+NVmgWAL5G3a2pO/vFp8/IwWD/FFUzPoK20WHvYD6
gWhAOg5jmdnK9urOqbhqOOJpnenOZ2aAypm0Iqu06Un6DMMF4T2LQm616tbhC++EMaKZJ1FOvoD0
kD1LikOnQEeAjMmtjAkxo3Jqh62khxwt1OC5CBH2L6Emuj1TdhQlrNHwLIw6LmhBAzYulk7kh57n
nAiOwjqoDMpg0jgclKA6BIqd2yPcbJpEeek2+ng0jJj1m89pdAet0Cb6cuGNsy2r9wHnZbgrDJ2t
7fi2CEriTxz2nFOVkXdcOs4xGqqvMycG0Vn7knPqQn/W6IwduWNBocrpdV89h8cecmcKU80K7N1E
6vxZXVGBiHd77s1NErJ634YLiYaEokOqllSyatcD1FxHjDLRHsAOAMbJZlr0k/sxpqrNQxu0EoZ+
XTnhzxON0abZKnEcQxzX23B9Q880QNo2e7w4iIAJO3cicaIAsdCLDmZnS7y35k1PgtuTMcGET7n5
JATJGcktjOEyxk1FZ0LXr1+y2aRUChpKUQ2H+ewFxxlo5IXI/M/MeiUBt3CPmdU2zZ/4QDS8wQnM
BIZafs388Hw9Vy4B1/Wx2Hy7stPXVH5sJwyprgPliu8X2h7PxHOJ/gwyQZ58neBkhERxvHnwY23h
AMTkKsqFIvJCN5D0iyQVKxCjq3iPQcQTGB7biJbd9I4+UHwTIgD1ngkwfWiMKb3zmqL7tWAd4l8P
wbtn3b/33X4otvh8TK3DxKlEYZ6svn0RVcn6fd2FPMXtC6/P8cbGZUBPg1HAIgUIiNOgkf43edBN
SIf3QRVNLQBzP8Ayu061op7Jb161Y12QEro0MT5wdnC+B5j22Ama+E+3ks0KtTNr9u3TwqvtB9g8
yYJLyqexKpxJTd+/w/Mpk2NOoWyThTmwlRIT74fwriotdsiir2bx4KqE3su0anGkhbLdj8jg5owp
2QK++tabXZRXj4uKpUZHeo3cWU7iYFW0uK3rbSdTWS80+RRTulTlE0hLTbQFh3NF6zhTFbRHPqLp
UCoO3HhTDWMEvO18gj+n7NNOAIqHEEqGDZ+wCk1kdQ1YwPe+8Wn7H9tx7PPf6myu1YHHmt6LdPVU
5cCW+OP+SgoZA0yVqIVTeJArRa7kktqprmHQQk1UCEOxAX5F0HLGNuwrpozVFRvsQPTfvO/Py82w
CNftlGPwk2K/HCtXG1y0SWB89oEhlqWgOvF92//AQ3DbvaePzgpSQjw4wpzRwk9ZKIe/1cMiCL1+
12GWAUu34MAtm5b29ns4VZ34He2eBEytVXJOO5nuXUF+ngVMYOX/2k/jDGU6Bl90Qkej+YBtRE8M
Adbiiwv2JW0CVTTGoLdbaeURNxJvXSpLm/n0zMt9gMTjZACT+46vNrAzkeGzVUELkDYzn72TPyfd
VVglwhiMMHjDxCoU/ZKIJh0jZJu6s4cZuV9NyetD3RTpzkQ7dT5/SVutUkYANzpICFB/oUS0ogpW
Fa36KFiCyF0hva3p0tpN8aMV01S/F2my00fGvQ8Ofx86utDhnpN6E7wOo/UaTWfAptNEEpp7Vq72
DDgAIsdGOqUmRHFWWS3LT37he3oylEM0CFUKu4PMDlfWqBkpcI1FtWFKzrYA+E/Nn/ozjbr6GPDK
mdjwsZJ9ok7uesVX+7LsdQOIyZtWD/bZ8r0ZXEyP1/eInGaVKG56P7W1Y8BsO1bSa6tE16tumXRk
vkuq5gSSTHE+EYU+70hPWamOzKRb1zpeBsrjjyC2JZRd1bX7Yxq1m0Dh5xbw6y+UvoAV/v7wJgg2
qQWV4m7fqpEzJBstNjp9nqwnrZqcd7d+XwyCjJ9NE8s+Wznw7NEB6ezPneZh988rRgbRJyY3kSnC
0BWvObr1lt90G+PF1k+wXN2LVVzzZ852NnIx8XgM4VkWIfTMnNKGLUiflEadfl78sRo1x/66Rkjh
ddozCXX/xU+TxCs3+bAnx+DNj/uj6s+uKrwHQYaRba2T16jDB8GYICLG5wlTpQiVKMPfJLCIEIKZ
aaNQrHRCk9GSEY8q9tBgU+wYd6L8visVPYWlMpQAxJumPif5At75aGtLrupeu7K55DStaKkI/WSI
mpIlv0EOLt073ioxDRe2SOaBSeVyTj6pjFelgvhlSigoqCUew4lmZPY9A58uaA4lXARrC4GVwIeP
i1ZingyNkJYjnet1YQSvMi2x/sKIQB2eXd+hfhqkXR2QRq8Jg9i8JyfROihSj+Ozebh9XCaYub3V
LyICjp7cFbA61gDl5ST6vKjNbCTm5jd74prlEwiOUIHPHdrplMl/p1ifvRHQciDUndE9PRoyaZ5W
sBcii+g7jGg6CgLxIold0aCHcsm3L4xpIbct/JEa6ny3xfia7EdxPen2ojKHzMOTzwzMpSk44ca/
aQGRXs5F+KXkdjTSa+omLLR+qxNF6jZXu+3OeP1hgxIjZVqOqPJjC2dCHbTi+tuU1hRF4ys4fb5V
hSoBn36PEECJ2J+KLZHoDiIN3eUfVzPexvCuhvYpMP7ZgilOMNUXMVMdYHrjc/ZBjrJqAYga0JQ3
9FQdP1ui/40iC7Ex+AN63FoIfiMl5FstHGC60RvXm85qEIYqWxZaIceSxDMIYz+Uqfa5v7hInX+6
ikjpd7CjMp6wzQWf7nVshRS3oN0GpV2nN0bvivud8ZDlMHAN+vm77a8qCDq/HqJBsj2GKOWQsqqF
XRkO/o70tt2asIzTBDLmWP98fOBBh5JaqVvRcMS+gidEgK7rC9GuuzjzQJ5RfpbYBjXghZh7H3BG
iDylSkEVvTnVyhABxUYxksbEyATJPQx5xYLvxHTiD6rM85FSPK6Mc6jaIcigUJbJIE9cvuqFQpp3
Sp/PxaV70BOwSsByz7WbGRTkidSvtPJ+v7+h3S+oJN5S5Bg04nlzCUzvgaixguoy6kqzxMpipzbS
B6JR9FO5bXvtxe2xtrXwu04W5xssgRPvKQA8M/4M/qUMYly5ebR6G7PlguvHWQ6dNPqnDtq38iFQ
263GPkChlajoLNnHivkFQBhZsmP/YfGMRqju66qUzClGoJXvWUOsJMdNi3Aivol4zYZUGdScT+9T
Fa2e2EsNtuEpNNn1+B2zzqhXd7qGqoZPQfg7jOM/MkDEodDSAbwqub+tm84gijMyLgq/sl8WplxO
banH7SWVQBtx1J5TDF2p94Zde/8ChnsG8I+y8KrdE+DzvxR+rsoPt6SanU1w3E0QIfV/Se5Y5foO
eQhASCQp3c4NnqVldWSB3JtcNKTOYZDoOz/KmKWaMQ539rXsNoYRj7im70WnMb98UzEZBwo+vO3N
RsKUW2SZ+zblygQ5pxe8wTLEOfX8BOP8vvkf1+cfKNEcZLGsL1oKUffZgtdMjYNZS9IYH1EJe0sr
5w2Q/H/dQBuWyXeOt2REvruOZfo7e49g0bfR5aYvZu8NLCknswAvM2hLA93kquTsOacj331Oqr75
w8fFxLQbkiabQlHRVB3Z6AXvHcT0Mu6lYn2rWdVmcDxO6xiUtwERvHUUg3ka1ujhh/IcIPjvcFO+
ZFHfc00NzraG3QCE6dS11+hXvpSY+5pzVevKXWMuQ7jMb6CjWS7SgxvCFC/JU3Lbuh+osaio9XDl
6bFF2ajX1gdkeabspBXn7t/n5SFiEzkAUzSECxUQGmtRAC+4j/6NMZM1JEEHxlLEJ9G6YJ84GjOW
n1Pl8avHDVs2eXlydjEBX2dbLcPh89sJO4UpIj9otgazCVDWV05GqRZ09vV6FPWTn72ApmeJb5Oz
/9qwCn5XOOOUXFyTgDUTW0Nif8+/n/0DjcpJWA2PIqgt4i8UtSC5y6l0cO2MCqk7T/xgcFF+fRGC
XzmrKqGP6gHOd7PoqzFqdrQCs9W5MBXxaiCkHFWjzTz7DFsJxtDWXlNoJQ/dGd5h5riF3W9jYwb4
XL4b+aknbbqcKK7Xb+xl8fgLDE3tvpC6V+OBHMlUkW9JZ9T4smbWBhTiOOmUWoP7WUmMPgzfNxuT
J4VVJuFdfKmZSttKEM/NiOvyTZZArHivG23s1C2wSBr+DMHbQ25A+7Mz5S51SiJN6PyYToReixDa
IYvHGvMfA3/wprkFUpwQwkKfm9RHcVI/B2HZDwCo1Oa1ixw+TweVixtgLtaNXklc0XQv4+NGd/+3
3U0iZ4gXJ1zU2ZFheA8TTYB052a1FKkzFjAmuhY9GrPCs2cktXkszcJ910J/HsW2Hv8m5xbkgj+q
sykjA9HN1SHFx9cD4yUzf66wdOWYwFidf0/YvfR+N2sNuz+mK96+ngQGmDWV7KgMlUc292piiSDd
Yc3Smuno4RK/Z2iHF4S85TbZmSv+Ih/81keuGbzj3BdAtGg44SwBxDHvRu0ir1qGr96//MSSwEeW
7EWtPhdUoNvqhMtUTcElHIMQrsnQczEgDojiuUrE9UjzGVWmtYdC8Ouw9iBF6QpLc6noN/kV4AGO
X2IfKCZ3mpVDWUHFRPNuB74Cn92bfkmR7AkxgCI9V0e9FR+a+er84hovtChn+RfMeQ9Ws61OLJ0B
cXU1vL3SmteDB4CHhdaONz0+2D4/Yjhn/oABC1Ygy4Bu9EUpW/wFFaOaDFS6aaamDa2g9+orPJds
Uzw6sweg31DVJdTSxDbXU8A3nQvUb1+9McST24ObLCOjyqrJE+bAtq+zQQIVkLmduogIdWNhThfn
xwIbdhGpc4aScaUa4rJJu1LZEXT96M18XZan5zHWoh1ORkZpeVq7O6DRuSfxUI4mlO87LGfv5NdZ
ql/N02RBOYU4f4HqY1KhCrkuDd408o387pyquWyOCycjnyjahWvyHDn3imd2KX+TLsNEgm6Q/6E7
oKPnzhcFmKDsJwF8A1JXCZuA3nPVQwQMf48jYwhiwT0T/Mx82OjQKyps1SxrCsK92Zs3LO0uOx3L
C4bK3jXclIpGNbRdd33hqse5egPICtcd84Y+DV/9JtON5rz3/8SZ7Ll+o/+SiKNn1CwSYwhAsORz
bew6krdhI8bgrP/SYV7ya70n0N/KJYIGDFM02iilB5LIREdBj8HuBeAT8rbcIFYUSR6CFCIVS7PM
p3KqRErkShE4vZLQvHfjvMmpfAr2eWqoq3tvw2jhubtrPuJ6Jc0tEQWPuGbJWPUeKGv3nA5pYrTJ
sNFu63aQ5v1J3vgE7gujuXFQRKoZYw5awI9i0qD8+GSuItrrDmE/2mj5r/s47lYTgUvD4mNPuGYa
m9uHx4aGKhjFFJH1jHcu9wy1kw5y2uvZ19hISWCt58rkuNrUqVtdGGq5yur9v8+4q/AP0z21ErGe
+RWe4v7zIfGCwnNiTkKU8drXynqJbcqMNog0fcD6Hew8V9tTTVSRxFvzNpKRL5tO9QMMUFc3qHC4
d8ZAGLwdywZ12tWYAXNdYkNm+u6ddiOUQSN8OfmFcmEzx6nvxnVSoplF7/tFvR/QOQAAMZ8qHU3A
Y/cvzu0N9KEzi0oIgDVco/sZujiyTUE3RCRtQP+a7Ue26Cboe+kDZ3XX8ce2fk//+1C8kg4ib+EM
3EOFkmhmcd9lertD9L4VPVccvrTf0qBv32tHcyv9knQMVrIJq3LxtbAvsrc3agcSW4PZe7bilDXm
gl77L6rBzMu7z0x4d3i4KTXGS2sxKJ0k/88pHJuvgMwfT6ZkrIa74pjloOTA/LuIvaBUFcTAaS9m
nGf4wCAwEDDHiyq1oLr8FFn50DR4MbTzaMep5ffIWulHx+dbde+Blp2Rcu8xS9PPpsI23B28F563
5Ido8abLH8A0jWF1+47gUf7WAudrhyubTI8LK0ICe0OoAogFYGOt048sOSh5BDKDpFYb5xpMadzE
pyXFxZ3PS351OPL8iMkKMXhOOIO9I46iw9HPiNlTJhiG5Ji/CIY/urWFQn2pjHtQDblhE+mrvO/h
Dw+o3Y3frugbAngcEHhPps+3/D43awJlrotgoEnsOi+xKViqaSaBq0k/Ge1h13vG3kjkWHcnnVV9
rVeb37Zffhmib6KzDgxOsO4ENYb5Pw3/bU23BCXw47CWp8bcSaxqdqTeq3pHK0LToOllsdf3PMgu
EHLxXQC8FEvtRZ0rBGtv40VkJ/h+FO1rmq2Hbyfze3a+iCVjTAa6z0vhzg882tLYhwNFyaRRSoMq
SV3RXZRplGVHJD49JkfJWJdXKVqRWWJU2G1XvZxJgIDY+m/99uv15Vyam91XcasQUlEOZX1vmfZr
dr0Nm8EMEPjyKY0BQXXQpypN+S16LzKetVEmwXJVlvktKqTapYalZJeE+lUArDzMkHMBtv479UQT
B1bkpg1Z8SN9wB0ZkyHcW3InKtGVpCY0pHReLNw/L/3nsBFy69bNZ8ZHSysvRFKwjGSaaDUw2DJE
LB14qAwT3Sj4zyXUKdvyHLba8TRw8edrmnTvu3jSMtOk4bouCD+M3lwKmz8VDtk6Ax4TAEn48OFd
r2cCAFoMLGEeGInWTohP1AsDGEi9jjaI44+q5jqCqPz/iplD3PjwE8+6Bao6Cl4FBppDnzldTqQc
z+nrOrBkZ29BG9hwTl8jPef+Nl9qZccPw/HrllpMSV4dQKjhPdTHecaQTmoAmSrapGCjbO3djVMD
mQMiNVwBKRw7LgxeAxDkmpc0mOcTwtdwkinwGVOmvTZFrA0+z4VNM4OAgRGVVqQ4rjt5wfkYxWmw
2lfyc3blOQtq+zHf1YrFGuhmk6BuSAp0SugHKn6p37R0TohJv2mUgydu0bksYn9e1to9R0NtXjZ8
0iExMtOO1GTVImBY5WJQDY5+/kUCHK6tPpT9SHQmccAw2RnQPOK3D4iBKLTtt532rMPNjhUvum/K
DJoVs5Y0j6o7Tyx8RmliBWUgkIH0iMoEdgwGnniuEVw21/uoMytRsytphpQrCiVpcB9KqM5vxQ1q
uKV8+rFi/zV7BMtKTJiALb3l/VpG6oNTbHHcwv3AYkfhQKAq8THJ/3eqOt9EvDlEL8Nbo9CjWsLK
8Fp9Rec8JmtyRxweEfoatUrXZXOcfb0Ab7y4BKvAyVPTzqlmIwno+B6whh+6B8bU67PFlQbKXNn6
wFpTTGd0eXJUE6vL2v1Dweeiia4wfSJc26ruSdQUAG0FD7rgit2emPCpbmR/4aGk0Y8PaP67OJbP
ttTTkkt8i+xrmamo0JjFRlP7H8YbZ+k+98AIsUJ8HV/0HD7EPCoTMqmRKsb0hOscztdX9R2hHWnQ
sxqCIRjeDfECLkS+KkXoilsSVat7v0D6h6D9cKHgS7uToM9g8PbPfg+KoOiwMCTuDKsMQRFdoUqB
pYihfgw6iVik4c73Km9X2Zg7FUeRNcN7r2oo2RTJQn/7o/QC5hp8gTBAiDenPcRoME+7JXveNeG3
WihTfygrey6VqSnzrLtZqmqz12qPPB6vFJTY73RxKzPp0/1mR6KFRwHeQIp7XP89nS72Uv54jEQg
XQMy9cGRCEheGBdvC56JSDRCAXdoELySPxNqGnCVgy9mhq68+mc15ZU75j5zpg9S7v+W6phFg0EJ
HcuhavD2uFVC1zkmLxnynQHJuUChlq6lqX7Z9XgYD9NgZx5l886fmUBeunynZLS94ntjYgvFbCc4
nfD2RxBGCkdhppxS+PXAjbN4XBWU4BXQ8mcvuccLrF5h++SmROo/fUAD+RXAYkCxLFUjsSFeJ4fs
RND9lNGJRsVfj/IjQNKrQ91L9k3/SFbs8en6pMr9BBNfjBtkDJZq/fbC6VYdd84SsH2eAjcLPtyt
s59CyW4P8G95DgyfBBdf12dp80oQ4BKyr6cjxGlOTb837/sjm8HghL1g0xCl8vTfSIjgkVoONJ+r
Jo3y7KwrofL6nH8nTSbGZUX32Zi0ji2Y+wsmYBOHwevw1+lTto1U9lb+ONItmmUWnzgAFm3y8hfw
jOzP/5XyS7YKGzqxCFwX8tVvUp3PLAwm4KR7kLST3/7cinjswHS4/DhDCSjqmTz4uQf4+ynDV4/a
9j+U9QchZ9FgAQeky8xQWujpS3XHxi4NenfJ7zhLszxiFYrAozqYdYLHSxarpK9YY4GiZt0gg74M
bI+W9BZAb0DXQdojq1XeYDacanqjus41SmcpCY0Am6WKFV0jUHG2O8HOQMymuEfryJyvawSUoUOe
AJR/Z+mYEKaxnm+2/PTUZ0NZ0R05E2tJzwovzIwr5WVIaAM3WSVyJUFJt79AvdjP/9P5jtndOCVw
FRsEd0oX1Es7vu3tMn4QrJB3tHFQOLh0723mPUrM/+NNEnB5c6MdkSZ0fTMFnKZSQW+1bRh5oclG
IOdGsWwstG2+TpJrFB+4ub3xqO2IbRdkFXt+vGfZr3Zz1lN73RyO1aOMfewtmuRIATi9zFnXDH1C
TsE1MsXCGzaFqGhc9WqGECzClwPqTc9yN53OKjAnugo5gnzUgP7yZbht9D2N7CgNVLP/sSo0CbWC
lMDUz95lx4B+dNIAJYjb1NR6zQlx1BMag9eUXfmPkdEssbErngeVI+tOTv5gOIq5KS0tgDj5Mwwo
I8c3denooxMNM3o0qJSQ8Bxd4hNfpxXY/6Qhkvfj6zEkXymB4GDMNqAfUifikpT47LEpQDiBVAkP
zCfCviyV2jmW/n6OhUpOrYdJIZL4QG2FSJVohhhkWMst00unNfJ1xRO6kfBwDXCYWyb2V9SZ8ky7
yCeBRrPvMNlBqKcYYSDGYdvzO8lBEsoiiPGWl+XyFTloRuXftz55CLGjNEhPF2ZpjBtQzo5NmAeV
M6S1ka/qirKjpIznxUIeOFBZUBWe822kf9Otth2B1c+tNlyyetUWwi2ouuIM8aofbymh9haW0J08
od/SeSs5x9YtsRZEyhXbskoHSRqmqvQfA+eq2iZJunX94NVIzeHHt0v+l66nH6BpatWNfEyAyPbj
NSzQYEyjyg437w9Uq8+AsMh9EshQqXVgjiXxAYq3YP3rFdsIZCauRTlPe6GlzlbB47MEnlD+VGK5
b5VceZtKd/h+uwFCuwiQb30i17W4uAb1JRhh7Iwl/JiPoLx8cb+CmIvfug0emYpxxCX3M8CoRhqD
JhNGv6Zka9zuOBNh0Id7fxKhw/Gpli6SjgOYOkrIQAA4+cHMkx+CzVHPxDAMJiKzEV7JYGODv97I
WmHHVoKwsMuEZtynA/mteOfl23rRq5NBCeJiRSCpfp+1z15YCeJ5PZlBPqO31VK3Aw8YqqdK2O5I
CFrefkwFsUojmvgoHaA8QGNqLuYSQYDCUufCn6Jpmbn0k+lJky+L+PeOYEOktVgm5tMR6hmirzFg
+lJGUmgEtmcoyncbUxeBt+OTiZGYIanEwOKbNo/yoHPZh8+ZoROYCisOdreHm7p9As4XvVvgYWA6
pdYNjS+MhaqgxiJPGNtMM3jd3GFPH3SyWdfr/YxfnszNkBUrA00fTI5IwvZYrN26pKDBwduF3L9m
a1sQPqLUYm//HjmgyJ08bw6DMtiEu12K7205dAqTQbAzA2LWbmV6xAobV9giuggs80LC/yHwFk7N
DAutkzrtLkGn+Nw0E1KAVyMyWSTCvQiE/FT6A7kAqF/6olikVaP9DgJtSxu7KmIv8MlOJpe/Lqey
ULKlNV31K16UnXkoWixJsq8eKKdNAPA5rZ9+Ei/0HM0SfYtnL6+KMk4YK7LPVgzPg+c0nredlxKf
WqmeQ6Ym/Ryuwylzz4K010SkDiDq4QvjyKSSFcy0kLP+dd0U8ibgPaWrHuu7U1RomTIGz9BRYvu+
hgco3Q9Ei5yv5uSuq+blhMeEjsJAYbVkoAxIXAtfLDOnnZt4z4Gm2mGFYDr2rYAY4etE5DxMpeli
INv9HxRgMXrYzJ4q7N2QcMBPFWd+tIPsOaanS2RQw05smAvUa6R4M0VVh105o/975k03Q9iUW8Bo
Dpsc7H9J9gof9JgSzGhnEP1Cm0pQ7oUZvkb0EdspTDX0G5MJ/BRjV7bRoE04+vhLovsHXw/IZ8OJ
/JaK366QtC0tAr7/2TVECrsQji0+xtVxHbFKfKYeR1+IcE2CtzCSi4JSvtvyhTh9YSj4or+5WQEk
xGNp5x3Vbu0bngqrkySC1z+r8AtmRzd0iHydzq9BGEsizMhMyFueEhckirn4WT7NTrfAGygd830g
0ASTUmyIYNbvOeptPyRLmdIiovEHuvzteWdMb1IailJYw3J6KfRJJfjqu097F5CqSv3DVzUTzOFr
HnZjgam4cLlvzqTVOXVDnVjDySv0nrRQaFHRel1HgGto9agjJcFCBHv3WHJlTS1AHR86RxnokImb
IzroYrx7Irm9xudmm2zkOBLcwD/Wfi3UPUiICEL8pWNTB8j+P6nPiYo9rIrKM48U4ObXcIOSsYaP
PIbaAEtOTjaVkHPtxP3g8nhwbG1DA4LQJRxkumyNe2R37MNS1WF9kzVDjGbEYMO6/RLbM7g0XKTJ
PgPVcYbbcBOKsgSb2d2mWkBPTYFY9ZMKKHEbUWevdK4zIzWhfRH/nBsPFe3M55WjvZHF2YZRB7j9
ByMhB/ZKZlFmG/8vK3ACmDPocDBb1/7SwRllwvEbb++3ysVXiSsgFx3UlNiBi8IZJbuMqWLP7e7F
q3LXZJvmP0ug+23qsOFItdCTKklhIz9O1lgnpMlEM0YTsWd4gFwQEOPqgZkHXO0TZKsPDJBdTJOy
0gLzhmVPrX+VyOs7rzKmkhdrXShOTScENIFhX2I4KQ01AI1XgpOJE0eIWc/zSMSzlBiz5ijPDtHu
7+MN6mumBXuO5c0N9JLftFuH008YdXyVR4xs1uCtjkGLwEtXBHdw6zfEiSoilhBSOLXNzrXtX4g3
/M5Yp8wEtUY3W0QvwN4W6cIL5/pdZstz2bRD8PnyMoIrmCSW0nYdV3zNJ6VB0Baggt6z87kFjGzz
+03G6sGbYG2ULQYvOXxDPN9PWgYTS3o2XFjtrtmTm28XCWyQPPf8ee0imXg5uVcGZRu1OKFZ0inx
sDbVlWEXH0Yj8zoUCikmKsHxWyu4KVrDYu665x3A+SRtYZk8EqeaOgkHbchppl9mPTKW4ZNdRF56
c7ZknrmdGQl4M/Sku1xVQ2VHfmFRD9BGadC0ecIIz6gHI/HuEiyrgXKUKxcrMZCTawSD7LS0eu89
uX/iohYLcvYuBy4wgJV2WWkgq261uveKmZ9eXB2RmkzGiKVBHdhglpb0+P4jkIUQzTyOeY9WQjUb
fQGl0jXwyKwcryN5ImLJhXz/J0jmgo6FqhKM5dKleeLcxBd9vT4Grz54EIL4mc+6cnAJbKgQeio7
M8LPEaU6G1anSoGZMyBFNiy9fnhrvY9ISVSGq1qCdwkFtm0BMPehu2kQvWn60RZx5sx/cvg6Vz/E
9/JGXFX7jEy+GEwt+rcVBywNv9DpJ6z7BpTu1yQjvV0V3YNW+C0wjqPo+yubaULgnLTeuLzY/xHa
WtBAHPz3vu4CRJ10QcepTdsgFBqA4ZS3MEKFWwfu3yyMy1U/zoF0P81kVUXAIoon2QwNAAae47fh
a02+bIzj3o4E1tW7ZzLWQ+4rLNZV9FqBNydqJ88IOzgqY3j8Ke01IH8YHaneqmrx/AqJS8uapuv1
oKbcWz/bTEIupTNdHd9Ox+IBJgRi+bXCTRhFebSn2koSLWLzKMhSn5iXhjIcM3lLTOBpUQcLLsIs
AcPzfMi4liUHAi2XNa/DhbMskoL2QG5eNNIVhZQbAjreQtiZNOBXSyIP1oKCPtLw2nywEBt2VkDv
vhiizo5xzxTE1hBbkP8sfu9nIO0JcV+BQsuB628a+lavHudN1D3pgloD8Ae1739azHcVcyR82N9G
wbWvyHE0uPX0jN2ZVoQ9Q0mjo1bUBb0IdU15OckPhNTKFwI+o4u+tFtu9Q42scXWBJQU1GsO6TOP
97ptbyFvnGKufh6ktVBCiHj6fsQssT0NOGwFbMe88+p//K2QLtg9w3EtYOu0nZY4TvIf4gO8YgYt
r/Ev2+R1c3EAuPaPAnM7cq1OsgJV0iX9BGRMEwSsdSx0skHnRMIptoiLe4eGUNwDJg9Iy5zuUs+r
r9F1/tbyr7HXC2QeJjeeiqV86kfZhlhOxnD3QmszbmiJwcDzK3IvUCFLUQXKn0rTAS+iuGluaW5T
OXajYY030UK8ioql9+tu6NDO1yueyLQ0MVROsXUqKTjeTAv4NPKFz/6yb8/2DE46iQUpnb5kOKJq
tpzxfbL44ecid9Sn947MxcsB25IXvJGcjvSSCNofd0u+VBcXFP87Rv/EAHwwNN6qxnxRpTLspkEh
D+q7QqOO6Y+InP9xbwW/LVRaOHyI6/xreXneZodsM0r+cvy/8DCSHCHi8Zd62U59txQCJxCGx/qS
bJsi+RhTWrLHAcFBydVbkPfS43iAkRAgUFkqDFpOjiWu9/oedRQVCF2UPHmqcAloz7EqItFeYz6b
HCYL6+eoWVt57C6dIP9EJW+om8GU7XyxZHPV7PiWNshpmPVoNAYbCaWfTTgVfZ5nTuI+w6XMW9Bv
bG2cnU6rovOvhIsn/RLbKzXveyV5fQFBekuYDBwT6xttiAGEsHoMtA0Mwf0PZbxJAzynVDBQ23Q8
R2PPyv3pjie/VSlt653rC2kZ0P8VStBDK0IvbrB3Ha06hxlfCdl3MH31MOraab98Xk+khTb/ZeeY
MxdqGhCSOqDK9m+UKG1vu22J2Wg3lBuOKj/LwNCpsqmKceiEEhMjoCOLCE3d5PDyAeXbhT7fPH2O
gdf4/BBW8qwEAz0FttozPfijAZmrigUxbjdkaftpuy0p0JQyPG+3S/+AnXOkDl/rDcfGkOAdZmTS
atdgnfL+S/DBRqdJ6IAsdRbE3heEUtGT+bMfcMNgBMjwmuv1EbThpbwQhzw0hN4Jzw1VmcBr/mh1
DDOEsHHhxPCtT3ZF9tYb7Ne2Pl1lQ+PahPZwLtRo3npYvBZqw7n+2Qmde1gDZDZAYm9dVrtY83bx
RsvjyT1URziMsw+FTaeXo37ZvQ2oX6zZYRK1KaCMFFwrPvozXqV6/jVora3M3izh1EPSgY83JuOO
jD9tSHbnv3UkLzrwywH9vVKU/EWTAUyqhD9gULvrlLBgz7ML2itJ6mqPI60INZQ/N0GG9TZZYXTd
LOX5YDo9QBy6JbWwbzSj65cDInHe+aEhLTvrcQPp9LZ0Pu5J/hJuMZ51K6j7gqtkmuXY3DoN1E9u
m0PKA6Ta1PMuDfW69141qfbEYEtEwrZEu2rOl52Vj3AYe/Cmqgrr+EiGMzF3Z/OLtiZiIsLSbmC/
8MnxZ5DDHpEl8SArp3ma34AKx1IDrNpK6ujJzCAWZn20B7RIseQaAkrOsGUAXhC/fMofHmBSpshx
18w2Ru/0fYfKT+2OAKKGqmAYGux9aQMyCGyrnTq31/U5Kugg/PC1p8uiMYzmNQr7kBAo2PN/oJlv
oq8LgHBnO17vh4+Ud3w6MR36+qoMvpnxYqRdxc+oG8jbkrewufXE1A3gLgamo3PKFG4/olm8qX26
Ikn7jsLHKQZDaMTXbur/G6xnN7Ns2KMSPNrk/sSsmhVHcZ996GSU4idOjKeMe0nm6+xFDEzKYP0t
Ox/QJIaAtL1LPWzMY0sp53UBDnNVKt8eqwQAEocx5iQGBdcbK232wM0DaoIxPmZcCR0yDneyWA86
CdQ4ZScZCpdThxu3c8dmAVyiJ3PZXTx2omu1oyLHXTukAkyK07rpt5seTxTnVQkYMwr0vv5jxbKv
mEAylGHXMiARrY4eIC9/4uFC2QgVY/1ieh/W0AAxAHYauSlob7FyitXxNPA7trg2zHQbdwPsJl5U
8Jzd61GS92uSzkDX2QkHg4KHUARmhQO0BKuYVYnKgCJPAoOLJlqVuaWvlMi1Be5zV3Ke8zIDBs3w
ns3kakowfiHx0CYY/cCRL6mM1GisiaiEGdw48zcoM5a2Xw0z9jK0I0QxPiMUKz1RgsgNey8DGrni
cz9by2aUAxTTnZu58fnEotWiSocPEJHcqfokz6KkOC0EHf66u+T77X54D7u0m+MMc38ycjXO719T
BJrkCKO0XCY2zcOZLQhi9XxdYj5eZBJfqjNIG0n6qroVq7YKc2MW+S0qkiH3I0pJYvLAO4NY4ko2
XWHNxcLPC4y1WjI8J6alrG2feGshub8cQX0WryJoTXynnAHZh+vc+xIeDRv9M0EgvlCYMP6jTv47
M7V0Ml5F8PUvTvfHt6aEuRd8gvVqmDGvHMg5uYpB9IyaSWRAGRC6eqQTxSfAoHvSrS/Oaew8gvmS
pOFcFeuH2Og+cAD50AzbMfK29BOVl/JuljGXvWToXYCbBRPKhDvXeWxgvS7aKpHUeiywwizL9Cc5
0ns4+7goIHH3G1eRTLzdwZcQ8wvSOriQZM3KH48noel0DacJkqqflNzCUzSx/B8OUvcgIPRfCZ9Y
zsT6LlOY9N65JresgR2rAP5IHLWSNqCZHZMwReTsY8U0gmTu9AWZc9mScjnFFiNElmOXQOR6FlHW
9zC2Wkt5D5lGcA3Lp33nUzF6xxJ07zPoxXQNiXEQQvZ6liJiA9qtv6shG4GaVXqq3N/JAr+ha4eP
WZJm+C1tCJNHrvZjXw47tiK4Nzl79Oe/U+eyDZ4/enS59gP4+i+xVlik7egc89EsaUbccxkLniR3
6fDXvSWc+MZ0VzoDH4t8Cj6xNdOpya1HZyrihYk4zq+zfrcUpecS70pbg5R4KstiZ0DpdOtgKJam
A4/6evsGq4QJAKp9pWcIMCnR8jgcZYcXWSboSRsNNPQoSGrS7X24St6q0gHSirPEx4I9J02SG9Pa
nI3XzyWUPO+qqN0oGGl3b8RfGOyxOkHEoq4uoWX6RytE0LscXXJmVuzBK1kd6HxkHmvoyVfDcWgC
xgZdnzkpYEXFEzQj2JRgrky3l7sSkXayKOJygNKzlrNGUnx4s6u51bUVB80472Dsewy45hGV36P1
3WDfLDLLyb5jjoDf9g5PIyN8AINahkv6eH2P9o+dCtmdV5VB4DM0gsHZUPPrq2/ri2fl4pIBakNc
8WHa6m2ZAQM/aFP2x3AI276NIpKc0J2owhlxzRSniiGLI9CFtxu3hWStPq4jAJliPsQLVitz9URR
g0Tgaa1l84svUMRyF+jNzRgH7tnWePmNciwmr4yMAd6uTc59O59SElH80lEKY7ZAE5BGfvD49T3r
K1q7hFw5xWx/CKbF/KKUhcNv5SSyJgzFE+wMK29zvjYBbxZ8XDuv+AeNoil8zC/FXlTPTfsqaG7Z
UaAqV6ZdkNP/kCiAIhA7UfupLOUQWLdCLZbyt+gRYqG0aOkOWdN7DUvisiSajFhKIOpA1CRkzQzp
WMpb3e0i52TjmM+tWKXP2f6EH34f3OB/u0NinrlYIzbm2NtK5IXzMNgNYutRx+ocCFlxUk4dMLH0
YDTo6LtO2trTC3EhrkfURYCPiA6PLi1swTvEot2QnpQ5/b2bsXyuTPsRGB56SYVG1c8uiliNXZzj
LwHjD5q31JbjxDUb12st4TFCBo8EE+qBm5VUUwPvSw5VXE0e7SzqRBUC6XPe0fpjdFNd0LE5n3pq
7IGumhscT3BTkbJWU772CQ6GS6zY+OXvi3+AsJsXSq5daO6bl/C1CuNTw9xtldbY4a9QZI/5Bqyc
Cr2JOERz1hzcHtYO5VCh06je2KwObLvptVCeCUdTybk4TIs8b1TPhbZihUKyJT0z0/GzQlS8SIi1
bE1f73o6kNlY65ydO/TFizLYG/sqB183bVi+bPJgSpKA9zWLQ2Vk89TW4/MMeyvKwcJwthsLMGwB
asb9+aGcxtCRVfC7Odw4PSc8+ESHc/ScjLgiUG3mk2ReYploxG768Jj8DdmFFyFPlGRYuCj6fspb
QeXJ12O3Q8oeu7nt6RNiPphJUpSH5YiCSM6uX7yygfq0wsuDrs+jZJL8pqFHnJBb0mtAyTy2Ffte
92ZDt5px8TVj19IAUW8/BmH29dFYMKbll6ulcRsAiC2r9d3mtq7kcWWXirzeU5vu7wb9QA4Dm93j
8oJG8TwFEGl+Tk6j2LT0xKWm1tS9FE8DNkhtvynijyaI9FTFsZwpm0c+sAMme9PS6DtbMdA8ZMzA
Y1fWZ+sxKSsNE3bK/vW2bsXLYuGQo3VXiTd0UL1tCSq3zHPxnzH3Uoczld2VIw6kc9TwH6JvMoia
eS1GTggdtZPItE696irZsqo72T0LnDhB0d+wxn29dyGdVYaBQ2jyq1m0jinBcguvq0snVoVVBJ+1
CT4xbtQUp0da6easOF2H125NHMInR1wOR9QDuPEpdZbJ8LFrrqPwW2bCJQuycjKXZOzLdhGDRHpD
8x7WsvgbAQLvDntTdsPwEkXltABPDj29bfKe/rllM7kXRlqH+lZnShu15H0H0Eu8YN28luFbONuO
zQIRls8TNk34bEnYPF5YHMJy5aR8OK37emn4qpzJpc9fwAo014g+3EiKkOzR+IAuwk96j7w050sA
FPvaRyPHAuechdO9rMq7iAFflZFsvR1K434ZhbtPBDXPOf1BF1aqRfEoSY00ztXcXzxumbri7g2U
qz6vj7Clomn22vVWrxLCZyrJS4FyCqnF8cRIgPhPXvpd/uRGIBhmSNRXzWnptP5VWYEKbXEyyo2H
9E/xyiXetbJCv13hCq4NiChLFL4nV0QUJlAcOVsl32VTQ6cKZ3jqt0SSFMfx+zJtI7YOpGVcRgQA
xZoW0EeUP8Lfkligf1Dzqu3gmoBgAHm1EO6wbqN9Xtr79ppdzMuG9LusU7jTJE3QEAcii6IFQSLy
yMnlZUj3GdWhX7yF322mBJmxplkBHUSieM9huZkBcTuamtm2TvQHH4P//RCp0vs3P5dC5OBjLXQI
7MvrlYKkHUNUz1cIaDcHC1vX64pqDPS6+e+jOJNfZMzar+tTdE3R6KxN3nQYGpaermzbRYRzha0s
cW8MLaP2+P2e9RqeYQ7y08t9wwIg5SViGLCR7zXdrAxq2Bs1fvwDTj068hJkJS2QR65O8OsInkM7
o9v2IPISPHeDCAuoJ4FRYcPUAMXOykrlXhb9EEs5DySXcYhJ1nWd7zokL52UjzIH1zBZDcWdCaGO
JcM1HvXH5bhK6jxGCocfFolNuKrlK4hIAmQSi63wWyMZW70Qt1Y2Rxx/p+SpQ2liD4m1BecuGfUr
llA1eo4lcdq2MkvD0l5CIPSvjAbn+f0XLDS6TQpJhMYdtTHb6wNHIjmo8spdu1uLhG24TW8HN7nx
QD0m12d5iQLszNGHA3bJ+XnfBta6mRWcLdz3DQuRBCd4KQU1Rh30dFVQIQ6aaw2j5RASn1ZddB43
Ep7ybTI31d5omQWqvz465yIhy1+y6lxnF0ausjz7QHk3yjxTxsiYu0rKGIUnjVXGsN/8d8BEtUPc
yuRTxRG+jntZctCNL/FW4eg+Rh1NO8SZt989zZfqYsC7uY+d8FOlqPQpNC3xi1SaMTYhXn4O0ERf
lyhf3LqyGkWjeMPE62PTHWGOc//UAGeUjBnl7iVF+wZxU8Wj4B76GHzeODdUq+nB7blMudOXK00J
90T14otFN3xEwSoVNwuq2+Rr/SdKzOnF4a2SqBs+qNtk4CpRSuXzPas7lRjOy95LBg/iS001t3Zj
GSnslFt0e7VparZpraI6PgQUCu8aGKUfYPk7r57oAQ5HGN4hkHIX1mkpqQuGefyKbz3aICch3co8
1R6IDnSBvd0xjQkbCQJYkUfOVfcmFdqhVjSRYOfe9ZVWZYV+BQdgz5ZtaBefck1pkp6tr7qXYiAj
pR3n62rQNSZoQeZvhJj0SeUdmpN4N3S7fo/bBzjg+t6m1jLpIkAMiSztqU/nyCAmoshuuArxMcP+
h/IHWJ7I3gw2o43/vYHa0IlResYNybaPo2IzWEccvgvsxDqeksAVrZRxPFE6bj2X2vdwEx1RiV68
YTziAZm6+ldYklmc745+ds+4iroUicyMp8iABmJMkRmu18HXZGWLPMWM/lyEcIYs6bOX4wLFkgDL
bz+1857QoBEV1NSTDDlR7K1/7X3GJiaFJ4J89iSqu9QdhkeMum0Ny60tabdTz1RnejYSNdxWWxW6
CJd2b5Dut6ZEpQ4KkEwE1JvtGRzCnHrAjHyCni6IfEG+lmXU8/d0KSaQ2euq4vXw4ZNu+mTTIg1b
dqpBrthFqa0Z5T3shN8R0gqwizl9ZbA05/epITzmAZ+K6TAvEkMjzJpdBdN0Om1/XJw3juliOWgQ
8b362ZLeXDk/lRUw1SjPC6rzACzYYda0KQam92u+m08yyDAWOhCriM0r86/NuckcSJqkylkI4tOG
3YMiATlEJsXOQZ4tuC581wqx6ArBd82Kuzm9ELRjnjMamejD3Ls502sNNQ/RpztKCkGE1rYaJ+XO
Pz6bPlE6ft4bcTkpPwMZXwgfSCz3kcQsqYiGNFI7DAvm+4UnHj/GKehbUNemDs/usgIgWVSGmtTO
+q/aneqMZLdT2p2qjuXjYANQNYK0wkzbKep0naIiBEomU+vwdM9+51OahPpP2KWpX7szdXbSQuSD
09hu59E90dP77BxgT3wcnaXXhl7OqAuUQD89AG1jzJWRtztMQ0uYCZl8sLfIygIYdRm9sgVjDLbT
sZIRCnTZ4hCjv5V1t1gy0ngl/621TVlIXy0AsC/EqFUujR64dHeKGBnsNyO9L3/2648bZXeumBNQ
b3eYFiR4F/TJNCTCjWq7O06i/abXnN75xD+5K9CK1fQLwxukjuV/T5VTwO2iDS2AYnUDkgLIEtdX
F1g8WPLC79/QNQZvjlql28KtRPzVnyeF7d+RLqjOfhPvc7w4weefuOp6O3eAmVhx0oAA70pGYoCk
dL20yymhYyvc/0QvNWK/NY1R5i+uwncNo1FMBwgSynADTu+QTU19RBr+Y1eTI6BGI7ZPLEzayWuv
l1Me4ylqsjQ0A52hdcPeGH3UmzoXTTo5R0xfJQMrkl410GO4DCGAoPmb2eVrCXrpQKUQFMLYkMv7
F68g0+x7n57uu+2UEWk6CJ6hdlla0qEiH4IESWwuiLxnHdCWVZPrGnnpVjA8nWyNJNl3EOBml53w
HBD3HaJEOyXaYYT7ShZFgSnLrcVj+GJPuZ697DMSJEqCO+PM0147q90bmcXIya16+eQPsk5mJIQl
QTUPTX/Jc+OHWC0QgF+UNZzvQsBvhfXmR87MY0GAXfDUkt+Uab3384WmCfObtRevoXBohnSlgIYe
hrv3aDj4kiL194hc2PtvL6Ap5LwtnWDvOYUx+kwysVT24couZ38EhvEwN4uXEG5MDjGTwcHMKvAl
hvE1l4llh4Bi75bJhwRtF8i+L0xT2OEULRsyWfdda9jJhAWTgifVQKZOUzkdMdFSxaUQRricFjbq
NQJabE69/4Gs3rk/ZOEFbQZotvyZtrhqsHxLHnanHH0taZ/CyDanAl/tzuEEUSnEL96mGehMgsw0
XSl6sjwD5BbeoRqq+mxTJAOZkJG5IDH+QIIDq+V4e4n0KuILjS2wIRr8FZJJlDNKpiFADVxdzPm6
g9dewbgTPEmEJBw67xcWZF5LsedXVzXDj2Wc5GmvNirdbvfoX1wBN8+sE99G0Y5fC12Rpea+kyJE
2tVSMegpa3lOxgXDMjuWgi1xmxAcDMt4woyQ/U6wnw2mkEXo9VhhfGeplpWy3t4R4bodQR+Nd5ad
39ReGDtVHXmyRDPFLT5D2jp+f7j2JaHiOmJI24PNYVGZvxyR+AkAiKs0jr5O9qtkla9NI+p8KPl5
3uMHd+mYpRJEwfBvbjhDRkM6JczFXRufR3uStpnWH+nK3Kq6Gw/uM+rFVmlPZ+d8l/dDB3r/zVQs
gSwzTFMHjKOGhYAF4r+XnvfyIWDD6TCCt6FbgPB13xs6aDH6vB0LWqbIwBXpbFDQHpU4AmJ4FfWQ
CBNlvJ8I3jy3gAZQ9Sx12v6UDtGHONGzG9dbZEPffoYdMjD3qvz8QW91RRvRbSNp6pzohRsFIFVe
/HUGklpvJ2eRFcLW8D16MFN4cwAhJDg6k8nhgWyiexymb7mquUTBRUZ6fu/YzMO0Zt3h90kzcdiS
5mHz9Aovzch3DRc8M0U+tI7YhDyPsMxvHHAMz0EW1fjEQxS8qkq+E41/V5oK6SHCqYqFZgyHCrPr
ZCjYBN/mKXQi9n6Na0I22cf0C/JXVfb+1wdx+yVyGtEwp7/CI5QTTAJ5dXUsIls2iNdAAh/dBhoG
TNr6XDgzkTqckoW4yBJwJumXbWKmP1W0KHg79sQkhwtHTHfjjHJn5BgayoNMf6HwJsVXwZGU29Qh
vQ3S54z956avvCNLfs1md1TKKc9vztDRYL6ORU/RzUZ4YSfuddvcl9x+JDQHg6jhT3ZH9E108+5p
jfT49AMTYWy08sy7S0m42yM5sUTjhJywB6ttHxPqdrsvecRy7y0kchZmt63FnP6Bx8VbIES/TTWw
ODOZEgIOLFJ8gtfP5qTbWT8zOsCbSXtlcTcjqep+tBix8dewmWopSi48FzgEDPIg8vNuv3NAyIu+
IcBj8Ml+uBXTvkRi5yJHu4hGEyS24L47jDRp9JeRiSmG8iTXPFfTcYmqSsdjaadxqRPZNkYZM4xb
8UDFs5Rm6Qe2Boo8cywtP7MvXMRk+wyOj70h9+VmevZYuZ9g10r2xS+W+WcSHWrIPk+lqfbq1BU+
NQYsiKC1tJy3hDpyzmwX+mRwzXGHL/sMacvsfBlDWgB5m315FpFqz2nfWeFO97+9f/pnPZh8p99o
Cu9Q6QO6tTlKefajPVzf6gn416O+uZ/Hl0VIpDGJJL4AvxQjOIK/VRP+c9XKT+77ecDIpWNrBRDp
VITeL730/B5XzZk0uhcrhtaloIl6XdvfYMhRbLbToof940gKaTf0rvSAS07IOSp0yH0gZ7b+2THR
WPdRyTzmOsweOA3Bdb5O3fWpDwTjySRykGOws2LlChF4Q9C+3eyKC6iFigTXx5DDCR0HVblzJra1
/A1ub5RYdbiXNIdSvwLRk31gB0uOXY0LUn0HQQAJ9fk2OpLk9QzzW02NpOQFbnpUXkknszQ3eyPK
+zwaXPfWUDNMQElhm8g4YGes2UAtwE9yqMZMBC1lYXW1m+MJqvtJ19xHVaDX0RRAEcXCUMdGCmLI
bf/XtonydPg7Hw2zAuWm/G9Fcj2rKaPzbuHQgyeddaM4bOGdIGd8q5Ok3R+/Zu9G5HarqCmrN4FC
UmnGSFTcqRo1GbQ+pFx2CmyW1QxiwYc9q6S0sETAQfZcCDD0FKxEG1ARCewuA8X4OIN1RKbmgj3J
uQGYoEZP55NZOeHvbUQJBRqi+sZWALcazhxnG8L6ep3ESmC0acYkzo3Yu2S6DQM5yjFjz2dC1A5X
979NpBNbE8DBhvWV+4I7Q/OMaAIG4A8uWmwk4T5LMnG+hrg9uwCrmOevHrEzTHxF++Xnb9DZg7A5
Edjm1j9YIY8+LPSC6QNVRSSbf5scMai+OyTFcFRGlMCOFVk7cjLmG2kBtXkDS0X8ZQe/RUFkzwyD
ihl3qnYTdsFviPWBwqk21dD4COQA7hSzx6ZbdrjncnPRLmVsJe9jHgeXAscfw+zvoYIjO5h3qW5q
SUl+IufzZuyxu5wImPv13HNFs6dyAZS/yKfgaUulAemjfUDMBj/EDoDLup5UJV5PE2IuFQwgXkxR
FXkBNSGAG63bHQotWzJFDpTMIaDoQuxq6WZ7IZntmX5v+SztXukuAAHG3rvyty9CmZ7e3/XB5lUm
Aj/ClLwzXhykM3PH8ps55WOcaiStla7o4am7WSodcvRAz6BH8hQpxMs0VI3q9/hieu2//hBrHwyY
hNiG7iP41bcNshL9897W8UfDWMVaBpfH60OWLCXtFJrAD5a1JryvFY4kvy+iEpFtOv1MdPLDldGK
5Nd/29R8zYlW6tT7kA/ctfeCYuFG50jhuTRnegtJPAvcWOaSBIriMeuMIGfW5XzV50GbpDSaXW0O
9eVSZatxhcx3Sckf+3Fi1+6lHI6kkXLAY6/hls0tqpySXKB3Iy58RlkQp1rWR87C0dB37SwiNOcC
ESqrlrFatyxit7/va3n2yJdV9newGeAzOAmQZ8oDjp9euClCURjk3o8lP149qRQbHb5iuKHLZXVt
O39XSHedJIX2c33KyddZYT7TFg8vnrRcnpaeDfQr/eulOjmr64DsvD7IcMuM0yHyjD6MIE8UAUjI
y06bQwvKf/toDhkXe7N1o12p9UXmOvDLUj4SAvq+a6Ikst8rCQyvkUGJUTRWaLx/tdzMt6wCJyDL
iO21rGJshL1TyNyI90ehAKNj4ey4H/noIAROdTdAgAQI78ykv+LsNJYIDCby8SM9BC+uF7EpFX7P
iheq9QxdJ3Vm40mMhIEJZBT9lpuQT162jfCY+3+nu3xE8E9rsR2+oVdnhgPeCKWu6ziG1oAIsbcG
8YKR+cZiYcp8hmmU29jrC6Qikz73PIlJs0DGITDn6OqCaOQEXTdOjTs4wgUTvEFpRfdtKiFwwZfJ
uXTYtbUBfvsafhRdzNee2kXKjeUHNNfqPUkq+M4d7xg1BS2geZJO4U8f62OTIG4R9jrV0Jx8Ahv4
GsoWEqLnhGtMJ1mmX4xIoC2lKK7yJS9KRfw4sIOMbtP3fVQKCG3WymP7NK/SxnvaEjVO9CdqWr48
oJN4/jHkpO3COlO04HAV25GiDYJ02Xql/+IF4J88UlPRe/eNb3MsSnOb9cy2wrHL0hIZyRyicuQY
giQSleluChmNUEkL2aZufkvE5sAqjJGg3pJSn3XuCWvrVavKIydts5TqldyRTRhyPi0A5vd9hs72
scZNtvcc10mOcKDzgb1H5N7o8Gxhhs/p9M+sfLvJH6g9EZtR/ljwUJ4vAHm5TTX8en6dVMvxXESs
wFiP2Sjez7kWnCjb/2755URDkpO5I9pmzIMOIMrCWJ3RYfZGJrcxkSGMe9Q3z5zCZNPSby4EvygB
4YTTsUSVvR1cMDHuHsbowSqVBRJH+vtO9c/G1vnuiSGI/61izjMkAWJMsGIRJsHZoXHp/C/Axbmq
B4ugHTE1Av8oAxTVHx+2fkaFNEfsmQ9xAwQ68ftMIFVawxAjflXKE8kXXeAX+XLJt0lZfNuHPYOa
+qKGUAHYMiIQKVptfzoqgjaEgaahdK2ndETJq0QOOG9t+1BT78a3S2OvaPOYtlT/glVxMcr3Xo+O
49LUK1gA79WuX3SOF/ky14af7w1n5IILpVzAu6cW3zhn8XC4jCYWOqsvrNmtyk/05ddIGrCK6PCQ
fW80blS4usVNxIdl76Lx33i1FoC1YkGnP0iYkxhxKKBkn5BUpv/oAANr1CWlE1873m1LBfTjOxDF
AmwtiJegIdbS5AT+A9lnAStLptc349AXLDHnZYABUB0e6B5i7uOOBWiL3qKitBStcMagNSiYWaPV
qwToG8Sk48X2Alf9B3wd7B1gG/N6LVcMQBQGqwgkXt4vRpkZvV2HQ8FsTqdOKlybaw1adMsU8cHx
9YZOTzQKLYiJu88jHLH/l04FEXHXXH21kWT4hGyCisoZZH40xGxnyW8JLIMj7mG1iWCuyYapBzwN
GaITm8X8kaUmQqi0Yj3Y04RYtQJlcr14hNuj5xP/AFk2o1o1NzT6pgb1Wm2EWhryL/IQNABsGBSo
ykqDaD70Us5UMyNOynYRSUgyqEh1afA5S4dBJN6XmREJcfnSxBIBt1xRBR6RTOzNr0Of9W1XNSDy
2EMcfzbhrwewQ92o9VqJ6k6pFUsjM+Qr9rmtrhughmmGPVD67L8r7tdFH3rbaCjsNVzxy/UCeUgg
YdXKT/+tRFkX/QNb9yKtJjTgcr8cc78Uz9IHghcwwqqhVoKdcTg0og4QDOmQbg8Aj0C0eQSCWN8x
G4gWppGMM6+D82yHL5rnEwBmUxDe+ak9X7sbJrQdBN/qgFJxiqrLUv2nNLu6eQdRui8j+Q0f7eeG
7E9sYU/WmIy/MFSRSe7JNolZqQP6/aUpA6OR3UpRRdB+ozJSJ9DAl9+itKxTmse8ypwMWxFF45c5
DgiLVM7tC2VDuRIOmjXxTk4vDVyAm29gr25hJZKbAYZrGa7TjJjpoQ5tZcP5ONaP4r3V1zbzF1+/
UvqftA5Qd23rjY2ivI4PNWvnpTNeqwXdxaZaWvpLg8GmXmq0Pb1y+/FyQuSlx8I54XlqF4MtY3em
Xt8IVZfdWk9PXAqG7oo87LQoNIeh51TtGAyvL49aDAi5SpJdHVYBf/pU9MT4sVNAEdDlJaN1Ii/f
SVgTeuovrgpDoYnNlEHwBq0lu3kmT+YEbF/vneRzJojDf8FKwDRC8Z5vj4mWSw5JXRDNDXVlQQj9
DykpvsM7AurGN4jAw73ELcUXpIMP31uqafkiYu1jowulaRBIEpWuPoPGoyqWsMrP7gVIdHzAzhlP
viYzqa10NA3yYx3Po0f1rTAiJ66uLhhc36IZfCB9Gf/UyQTB1LO3/PSSmGTMqdaXgPm4NdeWv0hW
TVGs/u+/IWjsasRxepQCBUZh5L2fQ3D4LGb77Z/zUNN2t2FTGyMStkCFMSmBrh9sx1IzVNkta31q
HIGnYGt4NTZ3vhHKDZNQnuYHzwpwpoQowm5H2V5uL6RHaMLczE3aUFT/fvg2igmkP7TFP6A2Zy9B
aboOXj3XsEAdfyuzRGQ/8Sn7fHvfg91OPvg1xHtnS2yv75C7LN5jdmbpe6VnNSqO0gOBEyCc+poe
gux38KlaF+mmHFGj4UOrxuCBmxVgoUXEGJkwwCGKwQieetoID0VWEafKmb1qBTU2/3rz0WuPhVGq
nuj/pDsuBYhehcJttF7fs3nvhm51YaESynZt1lTNCHkCDkn7H2e1kLtTh7G6+KT5U6ihXj3Q6eM1
o0nIgwjUhdJyW7+gyumq+UyZygLe8jCxT0B7wQ5s9uhdu2OniVz9KCw7JECtAhgiCSTMcuRruIzc
9CzS/7igoU2IAW6sA0E7dq8MJr6JOcqEnstZCxvP/eGIAePwxZHJ30yXUzYx+97UWEv6gNJzzyCR
JHN/IJi3J2Ejj5ZUn+zkAIjxncAh0Ws/xknCEF+P2P69URq5ONFap6+CSA86kaUmmWfUBEQ7TZeb
EpUzl8T71Of/qfCoxDOHavuZNGSEdd+WPrE8KAFzAnPfjVDGm9FdF5N9PEw0XzCXxkQs92ur3YQ9
720ZjIr+U6tabQd08iEfCRTIZ6Pq1HtVK7RQKUOeTO3TZKZnB1IjhYQYZxsjyJZ7aHKa3HU1fLb2
0I1ohMRSKCC2RmgdFqluGjcRlbQ1ugjuMlXSE3We1iSBIHWqIvr1BFd4Cwrp7fE11z4jxbTzH6ym
7TEZ+mi8ZP5ypQWtsUtkMn0AbcDLhAj/NlEGsvkA1InbQ4cYvK1KdesnfWd1vKFw0Jjx/SbFs9rk
sEDz63Qk/EGdRvZhWDKnSBDm0mCrRO0iDHrAlzOBWq0Aq1C6gViPSHIz3Ce6g4IK0ssr5cE62Q8x
hzlQeZ5NkFhClAFKTSAv7FAPGW3vab/rIshDHnwPzm+7EloXml8DmH9GLmr2mzoy2RbkXvABB4XZ
5YvJDPPS+6Pyw/H/dh+OYOmxM4hdCylwa4/rV8VEQy99kf0LHqXklG0FU3gNj85lVhItFY0HE4fw
UYzARS0JSqprtsYID7wmFt9D17WB+Y8ClqdvBk0L1WKLKDqV/4uDMJCZy1RYP1uUDurnr2D8RaIz
b94IoJIiXLmb8YH3SYAcUbLN7VvVC+snkIceUvGAD5CcPu7f2mSAmHggTuqrqnAEsoetiDKXmzER
Uug5Sxufw8x3sTGglLyECWfNPSIrKYsQNyPO26XqawA8n9SjgQ96mqWJ7Yy+kldTqe9xHm4+AyJn
GiTp1/ZSuMqV283FQPCoHicUIUuruW/4iS5luUj+0YniPp0TljZD+Px2id0UCH/T0Gu8RWycVBmG
qKw2NY/OajM6BWMD/Um1V80OKNaeBDEvucyOlogF6c9V1v3bi2SCyTLTCJDkjgUnpAASbm/lXlqF
A+mY03tZrrBJesJSWOE9zwq3To1cULH/ME08jL6xrkVbNdDdPDof3LXn/lSIjZWwVFN3CLGBbH0k
/dCy2SpeX280FeKMXTEYvzS6M8MTKeYbLlm6MiQYdwB28KwIj8VOZgQAlX51koqVwJozapv58HYS
UyBNRDWrkJ6psr6AZ92RuIT20c0V4VQQolxliCRHPH9zOWjCGK7JXx3JzuPvEQaQ5qJ/Jbr7NW0w
3zfIFqYkHdsMfoo06J8U7wnir7KewiaA8rRzsAyiPMpjJT2nN3cJrwj6d+GNVZEXFTATbYHI+Gku
1jxpQshm8XTksYJAAeQ+R10QKOsou4ohunve7Tzl5SXJo7DDZJUqnBfDq3I4D3NpaGNllLnxBO/X
iRNjXQJCu0M4NlQrgBMd2SsFJQeJMWIey8GKvzdDd6CJxoki5bg9C17RbJ4kLpaYFOTUyFw3uwYx
XdC+rd3b6PwvhzS7k5qqIAujgGXfyRZ+Ov5Y71LFvvWsAMHrpzLeLWE/i7RS4g9DhzEmtRhYdhXq
XPFuHUxS/pKJNPSSK/7acO6fBW5VlwOWUzKPmOmBORbwRi/4dhs+XYn+UcfnpC+o7KlMfFai84WL
WH6xPkQNv0uD2x/HZTe0vU76UbL3QxVZwXOzsiPPa7oHe3Wtf4Ml9vXfcmMp5ytf6zMGOVzAhJ1o
ujfTWLwd8ED9V/CfMNDLkMYxXEIqbuWZ7TiFrHZCiGj1L2GCeo7pAWWlvUgHfvJCB4sAlSA6I/0X
4IwoPpnPfGBV+kAT7ywe49NQ0oCp/Ddg/bOjrMQ7zyqmHXqPEytjGwvnbOvNmNpmdElBNHz0WxWB
Y+FIr2YO9uIiruB1KmsIcJBjWd5oiWkt44mefajOL60ydDzcCUvh19+wE5ZT2KoHNrfV5HEUQCDV
JlFzn7i7BWnJnUj1FSc8B2ZQ73jnrvUKZEbFFEqVXYf/pm7NMKZmf29qINrEwIbPImAf3wBv2noc
Zp5XGiGnY/LuouUFZsezBonJO2mYByQ3sqn9COs+/u3bDwJMRmCS3P9/jcbatk/ptmzIDtXKvshe
grPA0lRaUHxg7ZvZpSUDwd8Niv64CjINctSB/Q2RGpuwCr1+6lGOGkjU5vVfYWr5fga8ucfFToi2
rEo9jkGrTptofTqVunIJkYd6PEub+Aqfw4wGPsd/NKifCcZ48z75Zss9Bd8Yw/ZlvghJk7LVgq+M
TbdLvYZmLD3ep4oNIbEcUkBg0fjvTdbtKtPGNTc5c9AzQC0MHlz48mtqOOyU2alD3nVWpHX7odgF
pEZqF4AS+LvNS5Sapyi7K5dv3JuxiYMFvcIwLGhfme6zI4DmJ5KAFmiJLcQIMy8gMvk2oR70LH/c
3LQdv2fMzKAEwuFvd0fDscqdOThvUmwQrwGfoAlBziiEtoPoPyBCwC9emhBkEIFdTfmXUvgand6f
/99eOh0mRI22gWGvuFO4Iutk2SFybpzR+Wf3JEZJVdDjcwYJA+KpEZg12/CYjqc7XDj7GQysGI5e
ma16PR1P65Z7Q+l81eyfkQ/34kpYSjQ1Ct8r8kO22WJ4Glul7pGgMJp76gzSSmQLW4rlq2kOTP1v
cpeOYc97HuTV7csAl++0jR74CnU8rKXRqvzmSSvok38x8MNTzsae9SAQn2lXJSWBjFksK4Hg/7ig
JZg5o3qjOVoqViLj35MbgUG1H3Y0+fG9nAZTL+Z+LFU+/Cs+XeEnJxGanTDvdqYB8vPSzUWyvlwI
C4vnAdZphUNyJJVkYi4Nyoj1VPTsJyiCLT218V2XCG0NIFlCBXMi0Kvn7hMg1wSGJO/nYq7x97VV
4W70BCfXZcIgrD3FNspKzYKfUP3ulnfe3uxA79LA3PsiBvANdqTS3fxYDu4ZlpyLw158TVXN7WTH
XZzP1eP1tdILtbHXbzy/yNNXjqPkSikx3BIkDQJV6JyMN64JbpxculGJW4Y0ggd3TAFlY2Ik5wR9
BVPr2OaCAZC/Mu4pjt7BLyQEQaXT6hBHBi0ISgTH4fQTc5x7XhVvmBTaLLTvSrEzw3TYS7cgRQ9J
cQT/WtVA2uy09vVXg3yQwMpRuZ2CIsdPpOH95Ov9IOdBQv15UcHJGdLGdlNBMqhdf124hXiFM+z7
FqlZ2dYY/SV4oJkX/YJyXfqBi2WmthwYW3ttA0rfnq0w659uf+e0CbWOddUPxP3LFkQJ02KCV1oP
41buAnHqU+mgWwAM6j88z1x61x1WkNBwY73o5ZHnQvT9KzXquGuDLEm3kjRokCmvm+1cYDZfP8lf
bysBTnGpVEp0I16E8cTSy4qlWEZp+NgbWE4x2PUvgBzZUBgV7OjVc6gMJmiWDi0hqZl+sreRiTl0
xJnp7+nBN2FAfPdl8fS3Sw9id0EY3vndQ4HoGFjkibChJtp7G9fr4W5XRlXxMERXfpzrSZPzrETh
MfKq2mESrgUm6RYTDL6XYNGAlzXjc4cYigM6VMjwbapyBU5Q5wJOviLbLmTmnXU20KfcizzSk2xf
B9bm9Wa0jpFHHmU0zWAMJy3KM+HaNAXmOSeCy14+bprvsK/XEmZr6VFZN6cezq9LfzuaGaFcDGtf
G1gXfgQ2hmQrnNLYPE+xIVrXODCFn7F/J6Yev2ITPirzXoIQ7UErOcmcoxDUAEJvrPVpXteXUkkO
aFZJdgNBjlZtaKH7Ug0KG9HbuzGNfiaDa6O+xcvT+DceTyfOxI7oC3KgijRvxqGtM6frG2HDW6gH
AkiacOeH/+9yNZWsUIxeGtXCdica4u9TpU+A5p3a8viIq+CwiHhAHsKwykDr+ALmROAxJZd0r47e
0zS/6rn0LyGTCLZLY3O+ynnjOtjJIWYJ8MUizZo5fTlGZJe4M6ICwSXrBRm08CSzsX8TaHQPL4BD
ACbv+ehdXESCEicTnBEjv521JG2Z6eE4OOtaASaLjKvcsBat5J5Vx/OQGMxqkd5XpzGAioTtQwe9
w9368eur1H0u4Zt9OhzYkj2VUlpX6HuNV2DxXhPliyeocTu9bmdZtY2/NyHTUqxn5MufR+gzG190
g30WlWg+m2LvMu7T7uzaZhI6gdS6g2BVA9sA0oO2dxmx4wRvcZz7hAgEbhOKxnSti6rt1nb/3pvU
IKkhFwGcKMQjwVT4NaOo6a0vfKh6nKvhnt1I68VpV+hpzgk74dfHhJxVZZj1a0litVFQT+uixErP
3ZVUaFTXZajLHr+xvFmjHR/Wmfj/NR6+wevGCduvAMxvxcB6PD9dmSEWgmer1SUMMIB04VOhBnRW
h/I6E/RcN/Hdv3gnNhvXjhWWCSn6taBzr3j4ZSkwEyfH23zv+piwn0SvkA8vsxDAHxlTIebqdHZI
xx2dXmeS2G9gKcncxED6NaTJjq0CLKM9LusvNOn49JmmXNyC7G37Bp4HYqFGMUEEXf5cS8w+nrKG
lVQWY0mo2hFS+KX01T4aPdUGog4r8yzgyQ7H9r440Y/aWGIzKGceV3w/7vn258sMZd+KTsgEl+Zn
jwOEJQ3Lz7PuP+zj40IeUi2YVtLMZKS5rKD9LjJIHNkFZRNmmP8hlzZmuWnSGbqPQ/JuxxWIvXF7
2h5bLQGRkFk3MMJF+N8eueN2IKmIYQWKGEu7IweS2FoGADGQfQZZ2SzNt7KzECNmB0ivsytoF7hY
GZcd4waav1x4tgUlnHQNHay6nb+Kmg9yYFqfCBbJXi3HSb+pVXcCR4aXl6Y6ROu+KPApNM4BUX4g
kMDWMKMEupR0+YfTp7YLxx/z+QSqYDEYiRKbY/PEchzuYFFx/ZlXguAxiBhqlugRkv8OspQURcRL
RKxyJbLR8m0R+fzlHUZWpVTBW84dwiRvEZkKFHdS0wnG3oTTj3xvSRKspf2KYxiesUeXPLUtO/6e
JKm8u0DEmmxHwPr1KuvcTmDDzGMZt/8xbVW3OmsBE759cC0+6QnMR/JbC3bgV/i7xAZb+H5OAXF4
+yxMKTrtiN3bCKrpoloOI9O5CYQrUjeT+Rk4F1lEpJ7sjb53Y8G0Mcs9QW7tsg9dqdiu7PkDZXkt
eJDUYsSlQSqmNnm3kaX0/NlcNjd79JBVT1S5dDpBKZ+/xSgXIXzXFTvCEMbl6cbXd0mKCxYvCYtc
Kork61SCQPAv4FqTPhQ1Gz6UkaeJ3rrhZygwVF3+BoX/QgoWceh5dM8OXsEJ3Ch4myYGfJ7BvVGO
yDSw4TrQlVkcbm0RGp36N3/NZIyz4cmafXLDnWuDZR1qQaJqXKjLbO06JQ5zl6HBkVvXZE2ITa1N
8V9BvPmCielL3eJuOJGl7wyzRBwEizTe+Q2wyUBXL311LCTerDtsl8N5wF8beY31P7cHin6fV8sD
eO9ny9XHgPj0lG2B4zZDh1v2hDQBk2dwh9Cqs4GNFBz3AjArUCFXwSm3fn0ySjQbjLA5H6jaRPcU
FKLwj24FI94u85OxRPyTq6geCNcPNdwNdLYzdPYPuwGxtk+Z8YYP/tCscRmnljhdSXcv+D2v+u35
dLKFWM+l1vwN1QEqA8LWExcmVeYLga8CT5nIjW0Pn7qokFMhUnyjXsxk7MOGAhayOn3+gCH8UFnu
LQ2EK80PyGelCcVRhtAU+oWrgzDvlFNxlp3asFuXZU7iduATJtf5EBEK01nSoqsQcE+ML2q7TAyv
b1GKTa2KMkqRzlIKRRYEOkTOJ27VVgqlZCVpa7Bts3RCEq9v7zyI5fov04IzlkSnZPh1vkITddMd
03sZxVlW4OJ1meGtRi+MFo+Cdlckzb6j0vv20DlXL/o5McfZPeU5tN8YZpBfgxS2LdQalI3eD0wr
P2pV2bdPEtw+0dTL+ioiNUXBchtTyp01IGIV3gl6bKC/E+FDP/9Crr+halrP80c/wf7SdPUo2ROF
CaBcgzV7fEeUFvN1jT0IYoQ4t7XBjE5uaQfWPBKap7zuMiRpVjqKpeC/HgZCWLcuQVn0Ps1eeLcu
mSoX0PpddcwXGeGvVtCH3aRkQkFfnumO6hYsuJs2c/rw6S52RStmlX4CNHITDs6jvEDFJ0o7tdyK
1KeMUfs5oS6bGHBb3x9NB9J/qcwdxpPj88TDQTKaOvPfwsVT3IXRyC5VOyaGpWCMo9SFmtHk4RhV
NG92kLGAQ1j7g006jUxro/XANt9WSl+Ns1ggSE11UClaHaUgrkE6bEeY/stZTRP2iwzBTtcJ9HhF
tRGDrr+1+qgEC+H1EgQeuoo4LOCF/DPHcuxUiSvgvfkp4ZKz9m3Y7O06i6N/6HGrmFvuMAuBsyxr
RMhruWKcYPYEPHttrfW+1tmvn9pp+pGhTdZvHRj672BGGZ9VL9d7uVuHk4K0WfKVF5BiP8xor4nj
iz8nRu4TQkTiLWCXlLcS82T34e0E6KSyszlDnIK/e1/ne+c2v9b4TIHqSZVKLbMM9IsafpcrZV8J
97w3ud7HQLvSWOeN9jPWZgQ7bNuz3qgSS/za6iA444Qc4nxqn/9h69mBMFT7gRLKDwoIWE5cNPyR
VX4KBITeDoXsQZbCn0/oScAJj5kARo5ODB1HvWrSgcHFeIx7+JVrm5/6VlBJu0IdODYIFWX1nqWw
5aFg1qSXUaBOMxx7N6gaMNwVtw5XQO/QgCWpmlG2huuBeX3wTnxtIIyPyYLrjzehYwPAYUJ/PCGN
LuV6rgVGHM1uhSt/rPNSON7wL1LGep5RV07LFKs1vKsvDRaTdIunpb/nm2nUq077zDCuYUayx1id
yh3tRJk1JQlJzJxABR4lPlsZY62oOX0cb8uOyN3R7nsoAV7W5sXpfvL9p6oMRUiNkASM3jguMxed
hXfrP8yj7xO85Lytkd8JRCCc6FCIfal/86jop/rSFpRaXHpxmXY+En9uEE/i5FaYgehH9h6cDbiR
MQKbcIndBBm38SWWLcOg+Vyd9080zVfGONfq1x6xL/dAdBUpoMKCKu8OcGY8scroFO0DXRDmZZih
XhTJXBLi4ED4WnBi18oj4dw+LO1I/jorrpTE7Yq1uLuhzKZrwrbvR052/8iNPzqizw8YusgI8Si7
Pkt45uS14jX4sUgEVyJHIhtZg+zssZgoWJ7IGGf2lrr2YAS+7r9/rxTUjGmSfRr/psczmnS5KZUp
ogTAP5EivON9J0iN372s+7khOBzB8EndPpTuymQoxY1Oy0HXk1vzE7u2+AQspvDZXebZeOcaBPWn
c8j3hcsJLhHUgGUc2yMb6n4ChFgg2xO5bwEMmJhyJVJJJwHlti9L7GHqbGj4xAg4ipaf2+irvH7S
zyzc6QUDimycd359EF7AIG8fs7sBPO32QDjwFp8kF11jqs5HM0iDqureBklpVr/KlPyBlIUd2rHq
XGMJ3J6QrT6kCWnGxlBWvXl0+ZHNp0axaicNzVRqQ2U1oZKkEOgzdcWTVWqUGcQy7C495Gtl1b2+
EdKy5jrbIXo7robSYhHb5c/1V5qNRWmOiat2y6utF+QgnwCgh6Ke3qmK9uTFmkSh2hAl38Du1V58
iMfHY9V6GjwAJzYyI1iVPj4NPr3eCQfdVPd5oX6i6DewPQpKP5pK/bm+YnFCy7yjK2tRMevQbaQg
ScXrwztT2T/oOaRXQYqdm50MfVEEJ54PqlGyosVNDq8et4PF59xlrdl2FE2BWOo5B7Y3HermO/59
c+1WzfoINxjixHTM3PTh4+Y9gjS7DbnVlPE9hs9jRBDvnFdPDVzGYajeToSa2y4Nr7/kIqQOfqGj
aJMRxOvnWPZoguJZd0mJYjh6m15cYN1JWVSa0B/cWhxl6BV6Fb76QzVc7rl2ThQbbzagEqMwGHJH
Y+vzUFVPLYS370sxHwolWnQN27Ce3+lgfj07kezyTiX2m3KEy24/O/LyitvhxKeGVRLKUi+jmeot
JUpxqocoukGdT76wpEBxWhjQXnGq13Fp7M5Oyev56us1znK0l883mX/lEWRgSXegUju4ozQKc61o
8uLzOuWIRGFShqF/rDyw15QVMzstuYRhsHQu9xYHTcE4z9o+pcb7bfNqu+X9HhyeUoPdIM7t7CTx
zs6spF3Irj+UjZdJtb8NO/JihLLn1BIb9h0BsFD2ix/vzQbDd5wHURD6nlMzmOJDhmBKSlXxDt+s
9V9Ar+cR3aKlvo2w4Zk9Kfh3XlsOml2sQDLWDpVIqKacgbfTRSToDqAXbgeIyUlb90ChPxMVVkZW
aiHV0R12h1G5r+6my5Ar9PQxwDQomF//q0hhGvVCZkQd2VrwEoQg+orTpe03HIBPt//Mu3HJbGSZ
N3PQw0tO3HwSrkl4WzHVQWQxzkZgO325lwZObJN/xlqOhavdU74MnUsaXwNsAlHwZVg8WyA0UTed
9e3EVqkpjiwO0R6BSCy58XYbxmt474NQIDl9mfeRTGfoDzwuJQXWR65k9yeYBZRmnZsKV6S4rn5r
X5vytrQ/p5PsbusGk7YkQutvef1paWZwcuu4M4ZTCAWozrwvQs9229iBKw4B29Dy0MmbnNxmZ5OJ
tsaZiYSrj8Vevsr5kUFNyqLmfTbJwfL1oUp4LxrbyWpodNUusDZ2Y/bHzI4j2QpjRvkJZmRJczrx
rLAtBsEMiLTrQm9/gK05hjHc/sVfvw8rMuh6EuzLJto/KcpOKvj0Q9eRjLfvmU+BDxUauqsOwBBd
9CzCw3I9+lKZ7GT+PFnsOyfyboESAqRN/tyzwyviQ9Y1X/3cFPWEjSLEo2EI3d5trOCxF0u7osLT
a1v9N0wayOKFPu2yQbM6XynQJbed4LtKgconOm4LAYlSA8nEu+89WaUPjRuLuiNPFFQbQHsqwqNL
vdJmI635pLVJT8SU1h5Vpnp1ocnwTtCDX54iUdwMImVhDtOlm0NnjHpW3RSrflKKadgyIIoiVvON
xQGIUFZRtikao/cU+Ve4Wy4tunm349qMk71CASxUZJE8nBdwKXiw/B0IGrv+2t901DNthLiFnMk4
NYLSpODqK4UUBMOemwYAAk0xjjY+Ru5H3PvbmRIvfH40L68FtcAjHffga6m/LVfIAlWrqPiF344F
KZuGF92ivjORTxUyqCpmgArlAVN3DENWjUgls84jwPpp9+6WKypovKycoJDWnxe1yIZl57bJ/oq/
5SmlRwh9LjPReBFxPpVDOFLwgencR+cUFLflxI/qwrj5aomCvkQnpaIA0DhLIVl8NRpnyvzrYOvK
xLkKYX6t2TzUFV55VVvBfR5ws3sjS1vmGfSQy8boIU2zwiw9URO/bMWHQlb3OuhRN0nGgwtGN+cG
R1Oi1zUIYndCX4SCOG5Ed755yvjk3o5wkpaldPrkTyV2te5bDg2vupctsy8cRfzmF9Zpi7UhkH5e
NzxoAvGvTlJ3PKzIZ3U8kdosST1YAkq+nxN8rmIhGYaDSB+TwGnw2iql4FG38OMh8sfUbBoJYpcF
6ffqYXbpCoa8ur/MVwvGLf3rjyGKyZ2YkgQ7vmg1qmlLmixZ4z9UChwvdKcLpKIzQRpwyya/RNg4
ydb8Q7BvJvk+PP5F7dabyq+9Ptq0Y8U6F3PqmS69GXiXyG2NxRrPPrKwm58IJPBd+RiNyLnkczFU
nTK3hVz105fCrUw4w1kuK/1zZs9WrLz288qnA7ncNixkZZt5JOC6nzMuI69SFKnGVKBQ+EqnuFXH
Fsp26nN2Qef/YKX+makQ5Fxa9R3dTDc56gtfswhPSlrCsbbDUXBYFBXQksZXhAQk+PRIZ+1jvoRd
zC+DKX/p8JfhawAmQzRRNF2CFqF+VKrWl3GZy2xMzEIdNablsL7Iow3qcdoDZq1QD5wZVBBcQlhU
0d6pWi/lN3WVgTQevhf5PABTY+/vM2KfEWHt0lud4Kh0ttPioCK+JDRI8+4KXMrypv1A+ergbc5I
Iy15LM0V0wfCyVLASkQ9gdvbgst0ClVGuyGpZXyQL74SPLTfbMaNO8tt7oeWw6FWWk6V2IGKjtzT
dZKelr3ZaCkUz7WtpAI8IwTBVxT9lKbtp4P9luNhnLBZrHm8fNS9lcMUZs8sLI4RGDGWhXIabhas
Hc7tI5A0SCWvagPF3CsifBY4qvfVGSLI6WAUy8m2aAPkI8gukp7eUGM6QerU7k/R6nJVAcmkD4D3
yDZjlwopC2XjMqCMlE4GzV0oT82tp6KiIM8qa//Qw1Ol76zMwdY9WAZJZhuleLfci7FLAIy8bL6O
JssyRFiJysknw+YpatkuXNda2rw/C/Sb7Alnd1qfIPLXMbNnHZSitrZks20AFQjHo1ygyXMO5jrN
nQw9WgDKTSAgmVlHAGEvj9o/xsCMYimaGizpjVTMOvv0GCeyHovy2YqR3cibvZMgNmFlyfsNhN6t
U7aUOmiy9UeOiuIXnQGnQ6cd25IhmlPOAqp6lD2pdv8kCMV8OAoffgvQJCfCksavL+eSNeSBa63P
swnLr2+Cwuz14dxmYBt9BWk2ivO3hwhfDqV8+x5ukP7etXSF4bqvNFcYqr+HxkKlKypYssZiXMCM
duARgTXVecU01GdWeKY/mFwZHxVvp6HrZVybJoSjuMP5XPhPzO1wmhE7CJiWy2YUm5OYcTxkYeRP
NDlIW3jx068YjyhQ7t8putHQsnJE7ncE054Knho4QVZ5HmnQKk6uNHR09Y4P+tFnF1IVQEjwZ2Tk
DIBapPQNO9YeZsakmlGA8diknKlgDq5xJOqulJctiSj8D3EFB/ghrbCG3uFRgYbd1w4RfDRhLLYp
vOajcSzaq8CrRZpGczBXgDNB4Ygl8Zc74vrMUy0uHcO45UwTGj/2Pw9qIGbvsmIqovgv/6fKkERt
suqNp12z1WSmOVJpCOidTshyqny1gDVNRM4t1zcbay6UF2TW/szaITyZPrlI4pgYc+0QTQmALBUP
MV5s7CS5XjZXiTn0xWLKwZENBA4p8XsIbMMhcHWwIzHAgLqR0LSnmiEEKmDuYdEcXyJ5hsKs1u04
MIvvRUhtvBTrOc1wWKBvS0gTWgsAv7ZN20Vf8UMVHhy3ePWAAuRhEYhmtRzDxyiE6MW4TtNPprLl
4Ys3g8lDUf5Mq5BmeOO5HcL/n2tL75iegpYra0Dcdl1gP9W28jF4+HCgwocz4KmlLNTZHi7xTEhN
MA05lWoEBuoe/rfdaK2Yn9vBQBEcOyy7j+fP3HrWf2wNThRoeJt0DTg913/JVIXoSEQwwZPo3xPi
XS820EMGiyFtRs8kcggbSkEXd25wHZyhuAiqaNdlmMtSoRPLycYR1XHwYNZvMDex7sTVzkenaigW
4viCP4AwAQEOrV3aXomem+6Jp1e0niUrN2OKcNFJcF35ElvDN3CqO1j9vwYiQTxz4HgAfYWW+nBD
OQXGoKDTrYKz7BJ68CLG0Hk0zyBaomFB5Kizir9wu8FAAsUw7gm93TF0iTg1nrxD5qKR8V29IuYQ
zBCXGwDGs8mMgsbLOlovV0Vjsze2/o+5FWLJW3r0kedEkqZIiZotigCRNXeCA2yEtZMdk4XG1JLz
sLHd5Jh6hqCDSOGVwN82TJqtejPUSByiUm/eh8/bCMCZ8Fa0jzgTtGZmqQfnqOK3Q+QI6n0VUaDT
feTu+28YjlKfQGm8bu1UoYy16IRgB9RsWUCJUbrHAUoeRQTdqELDkxbbZxqJJi8ZxuTL1feLKl3O
T5GobheNsusPgE34kvfSJI3MLD9e1D8VtyPcY1RYtN+Y26vh+XXubampTddh+4wRtiONdpqvnIVm
kznUar0tLRwGtv4X1MJPlQEidS775o0dEVKqN86J8IbJJs0ICe/or+G6lCZiZwHhbLCQ4exZEw5p
76F/F1qvTAaBmUKLq+V/pnpbz2d0G9NsgRfzpYoNhwZKlqcslTPJsOVqfVDc2PyjzjjNB+iU4B+/
Y5WwlNbQwYL+MRGIQ9xXODvGx6LhhGE76l2U8ph3t4q2aHcv58A/mOMomuQX7XJmSh5twHNnlYqX
jfzEwSMvnSiuJ18JL6WODzcan5ZVKd9OYqY7nrpXHFeuC9PmHCqFy9eUdbWARAVJsfDviZA3kFgY
9GiPun7+FFcu7AbA5D8s8M1gm3UVJjgCu9CZy6AB5nbPEtexPVudVy97J77IX7cRXp/xN91Nm0Ks
tsy9jKTxov85oSlLPy3LxsvU2g6z2hT7FX/QbZrilxh7XAowSYsUxv2buq9L6NCeIAio+op8AdvN
2w8xtETtyeX6x+xw/ZXgymjeHTVlRrfsJm3qrwqyvvukKwuHFUJsAwHP/8L6dHOBrSqbMMwSDEcP
dNFWvt9N9WOgDyfJK1yncGAYpcjYTnCjFVf4qbnEEEixL4lBXhwHWZAe84+W/3vRZAKYVS4/dmWC
KeiKmmgupsDhvXBNDKsjiJq1UxFGCH4+fsu7EssGH07zUNlpRCu9E6rvyWYWAWm6q85fQRuLUqy0
qvMO0/L6cTBdNX3BZKxPBStnTYgZxfdFWif7RKlprUoJC2yCZ58VEkJ+SL05E8sG+gMd4r5lbqaI
V5Kvu5rsbn7uBrJzcQ4Glkqz/sLtRmwMeLRUGEvHG6xXkQKcoCWfkscybW8y4UpMzoEHlaG2o/A8
RF17rBP3FLdly1YUiHwDNmMb1V8X7KcvixgZV0pwtLmp7OQZbLREOcZ/Pgh5is9qKbFn4qdDtrsy
gzf4epmxFtBngBqJ4kmNFunfIFv74wyG0FvVIua4Oo6GPlPgO25NTdeEYPEKqeDNlRt+VO0QxwNL
VpB+l1B/4Vx+38voTLoyHvTYGZLypAdx15sqch/tAq972xNkXIIE054P/g3PDtI78r824GIBoN5t
H7iajGmgHWOPNYYyBePGlR8ikKRQ18rQfcQA7M6iv1zaiC+ZYEvcsd7w+5cEKaUHo/oUO8l8ibbh
84Kkke5uVl1TuwhOe8DhWhS66Xq4EnZgvmsr0lBRLjULgl/0CfL8ZI3zOcOJcduqGvRuIvN5X2Xb
8KukZm95njKYx7CfBqkUs/041u/HLdCPmjrKIQPt+D3wDJ0Xpc7ltNoc1/N+vArr6jgqXdWNpX+t
OgP0Kl0XuEq/8cLmo5lHKHW+B1+AxYryYV1S5LJYuNd4e4mw6q7gJFn1O6TOK42Djfnwvu4uDD+S
C6Y785YM8t+LOYhq/W8bCumQeQDkIl6vJrstPlxqnaU3PABaClm8Vf8XMgO0/PB1e7f+0v/WSz/Z
WzM0YdSm5b8tyvH5oOH81k24OPIClMC9j3pWIE/D1ISWR1Zzp28qdaBkPquhh4xtHsJGRzxeBOPv
BeO9vJv76K1wwaCEHUn8dqlKBzmj9hX3gw5yD/XqOOijD4TamSa6615KIqob/XWHrPlDEx/h6HEE
Th8hSTtPqDsJc2TVualap0qCpEu8GMdxdNhIP01jqeRFfKds9xGy7TEAYMlZR/R8K4euCgMniEmG
CTTkoaVOjGqbMaxpvc+6yOoo+GiWaE1mh15I2v5KuXhQSC/+A7I0QAkF6ZDpnLZxK1kKweb+Ns38
yd7tzz9T7lzHhB/kKrFBlqint9DwL6vKHC5uzgLHkorypeJGy3z3MVmZt3mMh80Kfwk/dz1yk7C3
ww+LD0VEdIFipo68RggJYgpYhdjvq35AXeHZkZQ9SGLOoczGl+1fXCvJP71eekoQqp2BVip7Jkn9
jf8vEBlzFrc3hcPAMCZcfeOR6yybRc1lYNrvyOvK2yXCx+EL3t8dOPCgubIVm3sHzlW+3McxGBJR
N1dbiTfT8Pb3pirzA6cCLPo83Zf7Jzj3rV/bBDIspgphTAQdSx/FMost5Ozhyihe869ibzL10tTv
5gmt90yrdCMUFtBuES+0vbGlsejBctUDderrVvYWkewgYU3YUQqlhl4kGfK6N908crIRxmGtWtIO
tNPcwE1iot9hAmeuQRBG/ijOIObUOPRvsVi63qcRVIcmOR9i0RxUDilDapecaDDEa0h6hEnayCWh
mJW/2FAd77lsfu0b2XXuEwOqowyTlJx2sejAbX+HkCqNBm4yaBfWDBPSteXx9Le3NaKgIWyEpjDA
dO+o31QEwpHWf8GiOAzFnoEujbagDrnjR8E2DfEYeOZQ4KZz7ytxYTRFeuHXmOIV7y2bntqCb4er
4eqc8Ts0stf8P+pvLIMRYmtUvdnKdTxLf5EIKa+C5FT4KVbQoj4B1B7938k0kK+mTBch/wS9VcxI
fJtMNsyyGf8lvQpfEAMW6Tz04baAm1+c315A3ecn9iALF4BlBHxLGtae7hC3HjQBSvlmi2HcZ26I
csMmCSuH7U4Qdm8nRNzbqEBqpxa9wbs7A1HwIAvTSm0nC7VVWPIxdxfb7oyagNslDHXfI38Q1mKb
ofi/oWw6UIvFlnl7InGSBwbjmDbpv6YS1ijDXswnapkwVTM/K67Do6PRnONWIeiJSDAUbt32WeH4
GMhcrUuszXzS6eFC8MoP9IQUww2QDh/oZTcXfNSFEOGO2tJku++wKHiSLhNamuKQJI1fRS0KT5jb
lE0EhvVSORsBKVuilqlGrQv1L8OqE4mpE+V3NStlFE4EAtlRpQDR8RcaTMokIOzOnRq9v2ljX2RF
6ee1mm5yYo3ADMqH9nT8RV23pZdM3ecVrM49wPc85lLr+Zmz90WmjyMcL03V9KBpnmmsT6HFORZc
/7HP6XRaq5UP3ecPSeyBWpwegNqt27UAAMYdVZqrC4u1zc62PHRRC98rfHysLKX8gVU3WH9lADBO
dec0q64hYDkAXS6rrRcEe48aWIMzMQVlfvs0FBLPwAbcuXU9xvkqe1UMnfqZj9eeHbXs6WAWkN9F
zHnru0abFX54E391PAKzYULvNnJJK5YAhDPt2JnpQwrAnAthbQ9MiaRU47Q75WvDzjxO7EQNC9r6
/ZDj/Buz+MGqYDZBbxL3e1Hh2612vY2xtB8mnQRcsVtWFSj2uhBipzu6yIIxkdZIipMsfoLjkPBz
Cs6wN1NwD9x5a54hBjsbIFo55Mu1kNSAkG5L9/PkqWEtGhSXgBg2WVFvxMAJAqw6dyRqpUyVy8dq
MAUqh3A1GLRPqh7J+d7Z4SJyZbR6VJZB+90mBnuP/PyY9AsWBryJ/ZgkqNvpqJRIQuiErhCt6bu1
c6ULgAl5gOR2G7uw8kI2A9o/sdzwTuKG2t/9Vui14/sQiQCT5ixtdTf8yPSChHsNsjMSlkmJXL2e
bhzuhje6oyGvAPCLBDsP+msnqprsJEdvyh7EY5XiBEowO8x14f9FAs3xLM5tClw159RnQMdt74WI
nWpblH7upcxN31KP2ZAZPzr8dNRKnsOkMx4uDGnrj+NEpIhyixiQmS0rd9dGjeuDS/2246q3oSmD
aynpO6fqtc/xXynm/gf3ZXECzc59tj4txFxuKuqbNgegZmQX92Q1yeCSG3A4qRWoVWuWp9tEWZ2O
dG9CuI7cEmpckzbX6nJhitKo7jJxRgjAKEfCpW+in1adLs1fPeHBz4Qiqvh7itd//5inOEuAMovR
TJYtUIdt/quxZancHPho+gDaPHIgDbqImg+N4YDQnc4haBs1ZP+3cTXZCWzVG8jJRvHeFFBSLUOz
XTl4rVgnSD+525IyWjeUcWu/AdQt/nA6j3klIx+WtntGEIg3OZ9jDdq5FiV7vFDRQdjyDVLobVuL
X1+rZ3Arfkpv8eWsjSVDDgMcWjWJUochmhcq8gkpokfOH/qQAO9KlZbh+BPaYa/3KyPIAT2zeeDm
SnORPR/wPUfMURmvUD/1ufjP1hWrxFbWHIpRGy0OCNJhQ5sLQfM7She42uLHqes+DpUZzdnT4Qpu
B4FV2zEC9nocJ8ADs+R9Ywc8kNRKCt2a64nPfux3Kz/tWuJMQ2J0VhsbeXaSmelyheMtkr3l89NW
omyOoqn6RhjQ5isO7aBu8BeqIaf+Cy8ixXz9komdoQaDkQ9SaJ/HPPsb5ZyYtjnq2z2x80y7niUE
umsbhPSDfTmEF49VwAr/oiu9XEY5dWTDWkj2r8jVsZ6ZFlJZMXBtpLKHJ+sntBz7tuwlWmSN+xW3
4u3esxdwjARbEiXHj1S0MXjFDA1Sikna3WG/6/4hfFPqY7Z+m23lzg3x7Tv+kY+XoXUF4/HqyUeY
zNEipVwb+nS1JXsyN+i2j8MbhmhYJ7yiK8L1jzUJj90xtE2rcX5lYfUzCL7UVYB4jqNd88yvbDvE
hciEKV7U+G1BDmXnBhjRz2EETE2OfOEzsOXsIzMnET3L8mOxoRxJ9N/bX3wdZMCGSci0utruEzSB
LwS+wQ13CzE0rJvCpZ0XczRhY1y+x7vao7K/sYS0bJiZfHc1gfPGHhXnVG3KBJVCMTTiXgxPh146
Zn5nhIuMsk28bTafw9QhZj8tfTJyJNepYaYItDqSDvU7bMlaJJgzZndiuNtsO1cTCeix9mVHzdqB
BfFVT5Eu2d1cquxyiO7i1mjJpyBuj46Bhz7Wqmc23KeXydNKaExQKRRwq33H0EsZ5qUxDHcvgoE0
fIE1NJDSQ5sYUdLWwd+HuEbDMv42FRORoLBPObE9uZGK4srBHwhHTipS/M12m4L4XZACiko/1YtT
7RWdpiUcIutzBvbAQeYHWnsBno8N3eFEorOlb7rPRu6m21EBh14Ue+7RL+7ok5CuvwRaCfSw8ubw
ksJH4aW/rb2Rs2zzbnvEK1Rjc8niUoOv9k0trD4sK5hgl4dxHYduuz1ewPnigv3P3BdtU3MINPAl
6u0u1s6noShqlcmf0PniWO3fpQ5WxmEqdDXHxZeGYBN4kS598gT3U4FrnoyACoBq6HxmJdIF1PmR
NvY+m72oABn1bGQt8DHhH7J2LvQTK9jEO9AiQhGP+TIoidFVMUlbF6l/SrUhclnuVBgL+jhnnSQP
ddBruKN0G/xChEFG6xObe8Rz1pITEBkPXxahRnobQAFOaD1u78xiILdbOXvfQa3k1uS0m9h7XWWC
URh0BCgA6ui+Hc8tqivft5IPeGSzV+KtYAZX8M+up8/b8DSfyAvWBZpsKNFmRaiBY6g9BtNzY7DD
uWdz7aZ5zwX3+Dj2z6FKdKAGgdgBP0lt2ezaZThtmo1T1lO1mco4TxL16RxUQZjV9GvdaRt3mgcy
0y1yoe8VMfpTHUN3qVIvf8Sd8AfQvM98ktHLoRTqT/R8+LQ2ETS04+mwPV7K2HtvgKpuPJFh5Xgy
ZtGsVfGHV3WA5XIiaWEVWzSNbRNeX+7AaOgbW0z5H4ZNmJX8mxkv8++a2Er9J5P6NrodFm3OUiPx
Yezd+1P1uSYZTEb/SbIVCRmmyeJoGElv795yNT1l0zOLHTrrzIny2AJKaAnqvW4d7kQ1rDBYs+10
+gI8vdVE7q/hHC+OPjtGH4x19l8/WWULC0nAj6dhNVvdSKQAv3L/36DJKiD6S6JOJQER0dlhQWnn
gbjAqoo2vDEPMWx8F/wdN21vQNiSJK3WZKyzfVC841h1dHfvmqBcILuQNwJqJCjs5j2C2cCRNBx7
w3VTkmVQsQNtafrCQTQ2qL3YvzQJfqh3Ef/nutMWQMb8mEkLRYBR8riwwEkrZrW70NUxr0BY5WYH
Zxh9WCsln91yP/pMAA39X07csFLHgBYwfaSpPPa5Vh5urMaUCuzljHJtAqStyqtEsb3unEz5SOLU
gMUbHRN3uC7KHl2wGukeKZ1Z/JyTjTvul8J/DetJnDWqwxSFOOD2fk9zSK4FBAH7TQmOT6yDE1Jx
a5llw29ccvaD57Y+OW91t9xhIgH5KTgcED09n/Rfqk6zc34bfrq/i0ZQhbfkSne0F6YDValJMiTK
/eb0xPx3sIA8yTCAdiUJcdeywGdHIWK/JLJAs2nkfs8prNtnwI9IPO//tZPL3ZYpNPdjyX65VzTD
w5l8/NNXM64Z9ZOvO43OscbLW84nxQqu3tUnL1/TDtJWV4wIepmOrMETGphyvYUap6j6N6BruVBb
q8ONVmxv5/5Zha+p34CntDLfbmVfThbjqbLRvKRiGSrj1SQGkasd36jauZ00QNDNTVGy5MxFhPXL
P1ixQvf0dW1C9GWMO1Oix3f+sB/25jzZ8o6CI7ryBE5NqTUEK62B5DZh+z9cVMn6frzp2Ggd89TX
9ql8MUbHUGgJ5YrpahV+MW2TQ0GI1mYJ5a1clgJlp40imy202lMB9kGWR4RfGS72ggP+CR9u1K3d
f4GJQyJ2m+Tf0d9am3BVuAYTkuTsVjzkgIyq/ch+Uoeww+/ftHRHW0LP4o/6fP6fww4HMEa7wHXl
/j1BcrZerGi3+pgaI0NPCUZbA+0vvOxMcNLSZWPi2Y0057/9589HEahP8uspY/uor/V7Je0QHat4
G09gpuJ/spdbQPPMpxoIYQtwjZHDNp3MlA+jgbZ2u4iErkUo5Sm8OQ5Q5A1SC7otJjY1mrOaG1Bj
WQRuQ8ZNEo+KQ6LgVCz51GKwA481SU54r15zitE2lrcf2e+WwnLvM2F8T90FhvfaAeCT6AFf+bQo
YgkW+H0nl/7U411Et8X/UZ3Y7G+YEUfUpnIKLxxdWWqy8luA6eGUSQnlJz6XfAB8N3dmZ+Z4U632
o6wWwpFt2E0QlmL5OkZUdMU8YY8oO0dpC1mNTK3lHhnp+rSQKGYOjAxfCKydwm7sXJ3wra0eFId1
cyJpWC1tgf6zuMZLivl4hWNR3wxppC7ApRTUw98JbmyI6CBqF92KC/Oe3P2R5m11d1722/drErNe
froO1mZ4lF8xZ0MRKmLIOjspTc65KyV05UcQdyRLxW737b8R3deLI4C0aFw/byeHpXotNdykLSD6
vGGWHtIJ56lKxQnOpSzdgDxc5WkPiGdWZ+m8CuxG0HAa+Uo6u+diJiXqvIsOiFel2didk/hAPQyo
u82xWZD6JuLeza2sMB9zohfIX7mma+MR8F5RB+rJ/ziFD20fJ18giV42pXaa7DCYQ5R2WiXCAZJp
8FVfrB8ArfxP/eaPSyg5+Q0zoH5TAWMxZO2wXg5AZLY5dI8QIuvUkCv2COsHUsZHM/A++HBl/iIO
3zO0yEBDOGnb+JYMx2dSyFrih7oub0Nn/7odP4FEPHGK1GMoDBko1MzS3KVlx81I3NFfJA/X26i0
MGklnByrE+70YSSaOhkE47tgGw2k+dsbFhiT4rJ8Mtc7ORYa4EWxRhOY1ybm5zSnHuNUhzsqpVf7
qyiLbteIGBK6gvVDcFExAZ5MuzVrHVKSzWg5/WhdXRtqqrkJZ15PPNJr8ER8m9gdgIey7L3iPfhM
OkLvPZCKbFSknM3qRFUIqYvOLJGblIfk3d6PVpp9549q34UEKRP3MkBFzeBFHsfSnABRDGjpDdZF
9CS3V9a8KFXX9veOyVj2rDLzyzOH9d1946geEB9wAgC2SK19IFVOkTue6XmyhNvptDOJh0OwGEA3
66waoM51zsflwZ49QbVB/JzdxkoW3YOk2MZ8GQ8cCxaVPYUg+FNiXnbmvnX7YGhBIdiHE+0cOo+o
1+6D0eW8y4aml0OwkBOGejORr1fdifI6tL2Y2tgxS839L8VqlYZAG5VmOfa1b9I1N+aFplxF3WXc
BPk+JFo613OAxR/6cB3tfZjDp2WMfjPNsUUVgNPbeubOrvqNIgxyKaTL422d7Yq7qc9qzyCepi8V
g3DZ1x3EtvuXSGoJUcSFMN7yhrOFwkjJ8a9D0WhY/4E2oiIhPrtEovmgDlECVNWJCcSPVoMWptyH
3IrW3xzZc17txonJC7Z4wGubH6PC1/QANjT0yw4K2EG6+mp8tKCLdl1v3rCuYLBNY2ilMGVPkfDG
jKXq/+uhEQYdChguKTQOm04OM3W412i3hmcPas5NFghOVuHs/MS+k76QclhRcs4Sq1szDbW+NXQc
AOTLgdoFwiaH+mfIW62BI5URKKwA4b963/aboJIfS9YwKVU/4Ua4hsgKua7J1tEtvF260VLQoamH
glc/+uplFOEjdODRCCKFXIeRCF/TMrVlIpnOclfO9dgotp/WNVAAU9CZpBmwssqZE6Bq5JEQAPTE
skqHJ4KR1FNzWTuEpX2tA/a8UmDqzjy5mlMjHPFi8Tgdm8EvOQmyW5bddO3ffjtl7Y6CoWYvLvPr
6Q8ZYc49flF7y6tfvoCzi8DX8Pgv2Rqi3lPSVDay/aRjkv7vO9oR43nLN8gd1gBxLlYS2oAHCBOy
rkzZplLyIa/lnwmVUQglZEC7q8F70q5xXQAiDOcHXr/bMbnVAaQc6GidSTQA8oFJUVpZLb4ezzlj
PwX3iEyJO5EFFmky6rWfnmxbXoZA/e41AtMBhLy+sReanRiQQyR8OHT5Grve4selhcCh95KZxKyF
0xE3jFudbIoQRzLSdCkzThb0lKm3vh8Nw14NGFfym4rnvdFa12JwbMpGFXFP/wHXpclz20NE7wLZ
8T1HwQRoh3MpremBvvPU5DBlmKYv7tRixloUQd1/FCUfJZMyMh6Z2hv5a0BHfUtahOmfVKoCZvus
gNYmYtyVENI2o4+T5FthYO7LDTMSlgIJ9bKcY+GM3tsGfA9ZGm7IsR8Jq5T3j26fY5Dl0tQjKzEB
PBkMJMYcqo9M2xfSs2r6T438OEHKQRojDQh6/qQVM2mZK205p70lSj7gGwCTxzBr56tkuPnxapf0
qQLVC3En74THuFzL5FcwUcu1yM3XLIIaM2hf4iiUGN9HSm4aYxsvjUgazXJQ4OodXeI1KWA/z90o
2/D8bl2xtvifvcM5u51oh4I2jAcbV+PbFku3RVxsna9WHRMUDtCs19fjVX5oXs1etkSoREU13nM2
7+fX8n1z3BYjzBqCYX7mQWuw0OKp4FMTD1BNdzNQL+jMqF3Og0asFCJqXiBGkfaOGZK14PzuBCQc
n2NsbHucLOqnknyVh4GSAd/s2c4kCFeSWQS7Rk3ZMKVwptqDoYbQ7M4858wIsKCgkg1+FLTaE5sh
Ua5NlZOs66YgPRd4JE8zOGw4H5ndru0u9CM2W6cv+DL31rjHAmz137XKTtkHu/tX/vXwSO1x1HW0
3ts5OqJZHskCRekhUyHrREp/56j6pOubyNCicedlYbYZA0DPhljkJCg1mLJFYCyY70hKCjH+cO9l
Sjyn8FCoSm4cAYNYUv6MVBgcRt/k+RoA771NGXhCs75DLOuMtz2xRy5obzwX9D+UK6vMM6LTHSGx
0oiL3zNDpjHEhsGqoOG3H4I4zaDDgPxJz7bwJtOa20fqbmKIWoxI3fz20HbQBtX8vW60BbXVNFbu
M8U6OhLYFExXcWWRovMIOZ9rqI6520LrAvaD/Ryfgzhx2i9EJIqCh4tyPvLS7qSogMjpNz09whwo
Iu0KLkUkAqDeYKrD6xacc20t9UMMKBYFy7aEiUOS8dGeaGoy+WNXFgPGLkBrtg2bZH6+dLWat/5C
YL1lpFawIcio07uGNdPKWOB6pr/Lk6gehlVr4mmy2MHF7k+HQMdE4ipmqwiZk2pAfG/AC2RGxUbt
fZ76dK1U0u0iAg0sQfImzuOyDhGdBdCnicuDeZ9VXoD4Gun+C5EZEHr7S30E20HWHbfZQukyg0Vf
ToRDsTFELSVyWXWtGY/6uOXq87W0Y9Ee5Roosr2B75CXlaiWjQ6rznPISYFo3EDd6921fDBaMwd2
UJNXEE35ZRzoyCC+UZ9fOTlAxtdEOq39ljs4Hpw8upPOfT1Uyf+i8+y+QkStSg/jnylmQWfcjq3p
ukrfJ5X2Hajfs5u6riSYqObZPap7MCj/rCpgAkSWky+cZgs/7GEhOIjGCVLT8utRHTX2cCqRaq0s
Im1zCNp+BHjoL5zUYBFjp/c5xLy2mAZq5DkH78VFmw3rYLsuTebc23NcMkshNzc+pbKvbj/DeBT7
XW7p6WOClPwxzA5dUu5lSMYsoto1G3ePz0jC0g6sZV9Z+9lhR9sage9aNzIeB7Dr5G1XvfK9oBPY
x7DPOQcxHASzE9gimDmdQHIpf+E6qdEgMdS+rOEzvY3uOV0tW4KWssrBdG4+XYHnnxm+B6PzFCZF
+2bsYBiturDsE4zQ/2Ls6Dd/7/k+YTSiG53dw9QUctobbWm0Cr+QAHUcNtQnbyktLNiBHm13HSIf
jUvib9+JGvqOgpd8auq5PKjnY/AuIUxqgwEvWJPjpGzZqkiyi3V7Wdgr6uoASeQ9TF8lQjrVlhLi
KIYrAk9j0tLE2sJFzDjAUPlJaiF2txez9rXaDjj97HJ/ESzgHy1w7ful5QrhytD3cdvMOBr4SO7j
Gzrw1eCuzuzXGVY/QfObOgx0sH29uuSVjlQEYtMbrEPxuHvDa/57WOP/t6TpCf8N2c2wZOoNtvL+
7iz/iRQn+yfyDPnT+DAV0aHfp2GzeuGOLD2SOpO0KoTcU7qoRGlR0aiAM3c4nf+p2d+NGYaKRxC0
ZT/RmPN+0G5JZHQR4H2h5h2nsloQVGYlsDOBNYq3NGSb88aSciLP53oJ1jDjEAmc7E9xcT04pCL4
Rg2EN8eUgbLJsMtLIm43hhOoR966BNsVukEkuTe7hcUyR9F+rYZ7aSRRNjRIe+xKSEPrnFHNOgJ8
1KehvOiGUU4Jd4zbQjBeH4eBkhTK9zE7PsSZpWSx/WCvlDKAXvm4LNwBqP7p6BwkzUh3yS6jO1jr
YLxZnhitWm9zaLOmkD+36fsreEVPMuUUxoVa5uqptwJ7kGECBjfp6F0s+sl1IzJmv0Im+BdVfP4X
kP0tHc9cW0ZrRpkO6T0QXw3IssGV/zd5vrYLzVRAjaeny0j0+pdLMpowafvgu/2T9Y37/DAT7sfu
YeCm2bsJSHz5P22Pm8B0mc2Dh5u1QlkUTF+MTewfCYaRWGkzCWqDW2CfRn+QM8EMCE+qDKec55N7
e3HGl8c4gkp6TGLvPHHoCJqFjjMMcoarokDGLcU/zpqL51zp5+7EMNTqlZVXI1AZeOROydMfxEIk
APAsqXYmLaO8/fAGiNKJcoXDAHbAjpHigTyJJBEeTrtnvAxi9V9i0scMAd6NkNAiem5JQZVk8Z6W
WMTACVcJfVEBXO06fIThFzAl7xwLNOhOMdPqKUlefV/i0svx6Gt4SkvSFqv5wzvGKc1oGQ5a4fuH
n0fdfMMFzBKZlgbLqWaem9xukA50AKeI+LPYqv0luTavKz3YED5PMxolIrvhbCQ62+vC5jbKmb/g
oqc6anoh93rL3HYLBR+m96ePRC4TagYmUepwj2Ur+4JLo6+0FInAv3E+veCa2Ixt7feaK9zTQ8Jd
/u8T/5cWjfwwnUTaPE9C6KfalWUA+RBfgZZdWJ2Ng/nKtKvtItQdax3rWMZhUGIeFsEa7YE8RIsC
2lB4qiuQCQis2egbwjLVTMd1RhiYcERa9v2Cmir/gpXJvtfaXMO5TpphCX+580dceB6LBOzaJJls
9rIvqA2kn0mOEYjcouVd9wt+WXAhQJVr+LzujcJQBCJMM3JRo66yMoTsQ454EIpuqSvVTOH+EMeO
15VxW6QGe6SlXq59nE7zFr06ZaCxM7U5Ex17Rn8V/W9VPNTVUjFX/8Ty6GAQ5awgo2tVi1uxNnJo
8QPreA/d3TlEghyTV7U/xVETitG5xKyEWQN46Qwnw8tpm2vjdjT8hPjbrIqXH2NmTSqS6AnBYamC
I71s8mg5MeIFvCtdQDJ/6XL2fKx40DK6HEVomX7XCserWPMWnbAfwVhJ+wZddO+IF1ENMh4xBQZU
d/CC6xr4Jyhpk95AheIp0Y061zDupOWXpD0qLJZgWz1Cd/nC84v89huZ71qFZmVzKamL7KYOo3bx
pJUQtJNNNOX1Ezn+C/4Whi+tLx4kaTigw2j++e1JyWcjolrYmaB31+IGXmavD9C7ex6G7nKqsom9
uwIduf1mqoe4Vm0BTwJKBRDBh57YV30pX1+HyL3i+ThE5NU3EQ3XE961X6cXI8czlStSjcAbF/15
D0P+LMp96tkWRIczXVtN1cs+P5s5Ygzgqbhm0GxZVxWzpDJR6pWGpblAEeI6zTMeaecpP0fuL4I+
HWZV7RmSPFK6uChJsuAUScDcRhX3lI9x7OTQBuf6mU5AA16vClFpB5ulyuF3dwqL9hhDpFU7rGb/
K9PzaJFBfHwudux9PCsWZYOlMyZv3hVtt8fRrcvCEIUPjpcEiRPvWdWyfnDJwudI2vmbHrNIQw==
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw5a;
use gw5a.components.all;

entity Triple_Speed_Ethernet_MAC_Top is
port(
  rgmii_rxc :  in std_logic;
  rgmii_rx_ctl :  in std_logic;
  rgmii_rxd :  in std_logic_vector(3 downto 0);
  gtx_clk :  in std_logic;
  rgmii_txc :  out std_logic;
  rgmii_tx_ctl :  out std_logic;
  rgmii_txd :  out std_logic_vector(3 downto 0);
  speedis1000 :  in std_logic;
  speedis10 :  in std_logic;
  duplex_status :  in std_logic;
  rstn :  in std_logic;
  rx_mac_clk :  out std_logic;
  rx_mac_valid :  out std_logic;
  rx_mac_data :  out std_logic_vector(7 downto 0);
  rx_mac_last :  out std_logic;
  rx_mac_error :  out std_logic;
  rx_statistics_valid :  out std_logic;
  rx_statistics_vector :  out std_logic_vector(26 downto 0);
  tx_mac_clk :  out std_logic;
  tx_mac_valid :  in std_logic;
  tx_mac_data :  in std_logic_vector(7 downto 0);
  tx_mac_last :  in std_logic;
  tx_mac_error :  in std_logic;
  tx_mac_ready :  out std_logic;
  tx_collision :  out std_logic;
  tx_retransmit :  out std_logic;
  tx_statistics_valid :  out std_logic;
  tx_statistics_vector :  out std_logic_vector(28 downto 0);
  rx_fcs_fwd_ena :  in std_logic;
  rx_jumbo_ena :  in std_logic;
  rx_pause_req :  out std_logic;
  rx_pause_val :  out std_logic_vector(15 downto 0);
  tx_fcs_fwd_ena :  in std_logic;
  tx_ifg_delay_ena :  in std_logic;
  tx_ifg_delay :  in std_logic_vector(7 downto 0);
  tx_pause_req :  in std_logic;
  tx_pause_val :  in std_logic_vector(15 downto 0);
  tx_pause_source_addr :  in std_logic_vector(47 downto 0);
  clk :  in std_logic;
  miim_phyad :  in std_logic_vector(4 downto 0);
  miim_regad :  in std_logic_vector(4 downto 0);
  miim_wrdata :  in std_logic_vector(15 downto 0);
  miim_wren :  in std_logic;
  miim_rden :  in std_logic;
  miim_rddata :  out std_logic_vector(15 downto 0);
  miim_rddata_valid :  out std_logic;
  miim_busy :  out std_logic;
  mdc :  out std_logic;
  mdio_in :  in std_logic;
  mdio_out :  out std_logic;
  mdio_oen :  out std_logic);
end Triple_Speed_Ethernet_MAC_Top;
architecture beh of Triple_Speed_Ethernet_MAC_Top is
  signal VCC_0 : std_logic ;
  signal GND_0 : std_logic ;
  signal NN : std_logic;
  signal NN_0 : std_logic;
  signal NN_1 : std_logic;
  signal NN_2 : std_logic;
  signal NN_3 : std_logic;
component \~triple_speed_mac.Triple_Speed_Ethernet_MAC_Top\
port(
  rgmii_rxc: in std_logic;
  VCC_0: in std_logic;
  duplex_status: in std_logic;
  rx_jumbo_ena: in std_logic;
  rx_fcs_fwd_ena: in std_logic;
  GND_0: in std_logic;
  gtx_clk: in std_logic;
  tx_pause_req: in std_logic;
  tx_ifg_delay_ena: in std_logic;
  tx_fcs_fwd_ena: in std_logic;
  tx_mac_valid: in std_logic;
  tx_mac_error: in std_logic;
  tx_mac_last: in std_logic;
  clk: in std_logic;
  miim_wren: in std_logic;
  miim_rden: in std_logic;
  mdio_in: in std_logic;
  rgmii_rx_ctl: in std_logic;
  speedis1000: in std_logic;
  rstn: in std_logic;
  speedis10: in std_logic;
  tx_pause_source_addr : in std_logic_vector(47 downto 0);
  tx_pause_val : in std_logic_vector(15 downto 0);
  tx_ifg_delay : in std_logic_vector(7 downto 0);
  tx_mac_data : in std_logic_vector(7 downto 0);
  miim_phyad : in std_logic_vector(4 downto 0);
  miim_regad : in std_logic_vector(4 downto 0);
  miim_wrdata : in std_logic_vector(15 downto 0);
  rgmii_rxd : in std_logic_vector(3 downto 0);
  rx_mac_valid: out std_logic;
  rx_mac_last: out std_logic;
  rx_mac_error: out std_logic;
  rx_statistics_valid: out std_logic;
  rx_pause_req: out std_logic;
  tx_mac_ready: out std_logic;
  tx_collision: out std_logic;
  tx_retransmit: out std_logic;
  tx_statistics_valid: out std_logic;
  mdio_oen: out std_logic;
  miim_rddata_valid: out std_logic;
  miim_busy: out std_logic;
  mdc: out std_logic;
  mdio_out: out std_logic;
  rgmii_tx_ctl: out std_logic;
  rgmii_txc: out std_logic;
  rx_mac_data : out std_logic_vector(7 downto 0);
  rx_statistics_vector_0 : out std_logic;
  rx_statistics_vector_1 : out std_logic;
  rx_statistics_vector_2 : out std_logic;
  rx_statistics_vector_3 : out std_logic;
  rx_statistics_vector_4 : out std_logic;
  rx_statistics_vector_6 : out std_logic;
  rx_statistics_vector_7 : out std_logic;
  rx_statistics_vector_8 : out std_logic;
  rx_statistics_vector_9 : out std_logic;
  rx_statistics_vector_10 : out std_logic;
  rx_statistics_vector_11 : out std_logic;
  rx_statistics_vector_12 : out std_logic;
  rx_statistics_vector_13 : out std_logic;
  rx_statistics_vector_14 : out std_logic;
  rx_statistics_vector_15 : out std_logic;
  rx_statistics_vector_16 : out std_logic;
  rx_statistics_vector_17 : out std_logic;
  rx_statistics_vector_18 : out std_logic;
  rx_statistics_vector_19 : out std_logic;
  rx_statistics_vector_20 : out std_logic;
  rx_statistics_vector_21 : out std_logic;
  rx_statistics_vector_22 : out std_logic;
  rx_statistics_vector_23 : out std_logic;
  rx_statistics_vector_24 : out std_logic;
  rx_statistics_vector_25 : out std_logic;
  rx_statistics_vector_26 : out std_logic;
  rx_pause_val : out std_logic_vector(15 downto 0);
  tx_statistics_vector : out std_logic_vector(28 downto 0);
  miim_rddata : out std_logic_vector(15 downto 0);
  rgmii_txd : out std_logic_vector(3 downto 0));
end component;
begin
VCC_s11: VCC
port map (
  V => VCC_0);
GND_s12: GND
port map (
  G => GND_0);
GSR_4: GSR
port map (
  GSRI => VCC_0);
u_triple_speed_mac: \~triple_speed_mac.Triple_Speed_Ethernet_MAC_Top\
port map(
  rgmii_rxc => rgmii_rxc,
  VCC_0 => VCC_0,
  duplex_status => duplex_status,
  rx_jumbo_ena => rx_jumbo_ena,
  rx_fcs_fwd_ena => rx_fcs_fwd_ena,
  GND_0 => GND_0,
  gtx_clk => gtx_clk,
  tx_pause_req => tx_pause_req,
  tx_ifg_delay_ena => tx_ifg_delay_ena,
  tx_fcs_fwd_ena => tx_fcs_fwd_ena,
  tx_mac_valid => tx_mac_valid,
  tx_mac_error => tx_mac_error,
  tx_mac_last => tx_mac_last,
  clk => clk,
  miim_wren => miim_wren,
  miim_rden => miim_rden,
  mdio_in => mdio_in,
  rgmii_rx_ctl => rgmii_rx_ctl,
  speedis1000 => speedis1000,
  rstn => rstn,
  speedis10 => speedis10,
  tx_pause_source_addr(47 downto 0) => tx_pause_source_addr(47 downto 0),
  tx_pause_val(15 downto 0) => tx_pause_val(15 downto 0),
  tx_ifg_delay(7 downto 0) => tx_ifg_delay(7 downto 0),
  tx_mac_data(7 downto 0) => tx_mac_data(7 downto 0),
  miim_phyad(4 downto 0) => miim_phyad(4 downto 0),
  miim_regad(4 downto 0) => miim_regad(4 downto 0),
  miim_wrdata(15 downto 0) => miim_wrdata(15 downto 0),
  rgmii_rxd(3 downto 0) => rgmii_rxd(3 downto 0),
  rx_mac_valid => rx_mac_valid,
  rx_mac_last => rx_mac_last,
  rx_mac_error => rx_mac_error,
  rx_statistics_valid => rx_statistics_valid,
  rx_pause_req => NN_0,
  tx_mac_ready => NN_2,
  tx_collision => NN_1,
  tx_retransmit => NN_3,
  tx_statistics_valid => tx_statistics_valid,
  mdio_oen => mdio_oen,
  miim_rddata_valid => miim_rddata_valid,
  miim_busy => miim_busy,
  mdc => NN,
  mdio_out => mdio_out,
  rgmii_tx_ctl => rgmii_tx_ctl,
  rgmii_txc => rgmii_txc,
  rx_mac_data(7 downto 0) => rx_mac_data(7 downto 0),
  rx_statistics_vector_0 => rx_statistics_vector(0),
  rx_statistics_vector_1 => rx_statistics_vector(1),
  rx_statistics_vector_2 => rx_statistics_vector(2),
  rx_statistics_vector_3 => rx_statistics_vector(3),
  rx_statistics_vector_4 => rx_statistics_vector(4),
  rx_statistics_vector_6 => rx_statistics_vector(6),
  rx_statistics_vector_7 => rx_statistics_vector(7),
  rx_statistics_vector_8 => rx_statistics_vector(8),
  rx_statistics_vector_9 => rx_statistics_vector(9),
  rx_statistics_vector_10 => rx_statistics_vector(10),
  rx_statistics_vector_11 => rx_statistics_vector(11),
  rx_statistics_vector_12 => rx_statistics_vector(12),
  rx_statistics_vector_13 => rx_statistics_vector(13),
  rx_statistics_vector_14 => rx_statistics_vector(14),
  rx_statistics_vector_15 => rx_statistics_vector(15),
  rx_statistics_vector_16 => rx_statistics_vector(16),
  rx_statistics_vector_17 => rx_statistics_vector(17),
  rx_statistics_vector_18 => rx_statistics_vector(18),
  rx_statistics_vector_19 => rx_statistics_vector(19),
  rx_statistics_vector_20 => rx_statistics_vector(20),
  rx_statistics_vector_21 => rx_statistics_vector(21),
  rx_statistics_vector_22 => rx_statistics_vector(22),
  rx_statistics_vector_23 => rx_statistics_vector(23),
  rx_statistics_vector_24 => rx_statistics_vector(24),
  rx_statistics_vector_25 => rx_statistics_vector(25),
  rx_statistics_vector_26 => rx_statistics_vector(26),
  rx_pause_val(15 downto 0) => rx_pause_val(15 downto 0),
  tx_statistics_vector(28 downto 0) => tx_statistics_vector(28 downto 0),
  miim_rddata(15 downto 0) => miim_rddata(15 downto 0),
  rgmii_txd(3 downto 0) => rgmii_txd(3 downto 0));
  rx_mac_clk <= rgmii_rxc;
  tx_mac_clk <= gtx_clk;
  mdc <= NN;
  rx_pause_req <= NN_0;
  rx_statistics_vector(5) <= NN_0;
  tx_collision <= NN_1;
  tx_mac_ready <= NN_2;
  tx_retransmit <= NN_3;
end beh;
