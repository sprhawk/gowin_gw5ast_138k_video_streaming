`define UART_MASTER_SYSCLK 5e+07
`define UART_BAUD_RATE 115200
`define EBR_BASED
