--
--Written by GowinSynthesis
--Tool Version "V1.9.11.02"
--Thu Aug 14 16:04:06 2025

--Source file index table:
--file0 "\/home/hongbo/.local/Gowin_V1.9.11.02_SP1_linux/IDE/ipcore/UARTMASTER/data/uart_master_top.v"
--file1 "\/home/hongbo/.local/Gowin_V1.9.11.02_SP1_linux/IDE/ipcore/UARTMASTER/data/uart_master_encrypt.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
SWdx6Xds8vAMF2p7oT1FD6ouM56KluVkI+Ik3c7cTQPHJAlQGrHPPEQr5t8PNWYhceFD2cdu1IsC
VAmGdhVH37NgHk5B+B40B7gXwYbX3jpwh5zCPwiew4Skjx4Q+mJ/vVPj8e+e1oBu/CS74Mfy4i5S
rjw0R/+1YGfUvpefUF/sFWuxRnMdLs9mZ+gvBpitwt5X45P7bnVHfj2TnU/iBs4fuB2k++WzUY/x
InG5JQpyNnLeKsuQQGzSdH+lVQx88nIsTTssVCfICYB3RQ+KoajlWcb9OnqHekGGLoa8HeA95dKU
qLjJ02/0MRLsDupWuGhgTfOyXjczVZA1TiEQfg==

`protect encoding=(enctype="base64", line_length=76, bytes=107712)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
92sODQBTNsr664AH0glW54DYPzzklVdU3Hk2/Z8xgB5jSJZcXPQs4bagjSDzlysnX9tTsUXVBPsz
SX/6RBhk5HDOrEixqAPIXuiR3CSSZVWqVZRY4exBfgwBBNH9XOVax+0ymr56fyDOOuZsh9InJUka
W33jA5f1Fbq59SuiX9lhE/ouiyi/7plC2OrA8+2fCCOx3T69r0ZUPRF5DzilMInH221L5hPPp/ho
krljh5NPzN1gQgaGTDWavE/boIddjCuHzQPZRQGhW7e7NKuKIgmiu00C4HxiNo7BwxGIg9jsKJ26
aoIPpzyZQK8++zJN3lSonm3VHys1vtxhmr7zrD7iXnNh5iHxK4jcxS8ohFK4qh5ApRgDqrdS9n24
GIbZda/G15Cd91A8MNgiDJkVm5U9RSoALV72N3Elo9ae+uvAtJztHT40jyXOFQHFeYg07qVJDx+A
4UJhF65l05fQS8RJ1hnmS4p/vv+WBmYvUqRBv8BufTrBx6+B4dhNIMsv9vD0b1OCk2AXOIpSP1G+
nwDSEJbkNNY7ty0LGq4I9JD0+ckzBo6AOyKsfbXYxXnbXYBhIAsEaT4R4BOFJxwfJfwQKoZjbL4b
JQHYQHIE/OXM1K7eRoyQvf7CscvQeuJfIDz3E6dHEjcAvLCNpYTGW2rzo7xO9mxyfl/SN2vzL7hL
YAngnyUbEK/Rtb1Y9mcLI4d0NX6KQ0HA965bHg9d2UHt3sZbRr3vxR11BUQkOAPza2Lkj8nIgLpL
2BuDxepiFx24h/R6sZQ0P78oLqZ2fOjKQVuq2AgGABrpcP08SsluBDqaVM5F/dprrIXgStHoYWkd
JYko9NOLAlnE8KzEJphHwatYzfllwzJbwHTE4MDxLDMRfgKpF5sNL5uew9dgkxwcKnvEueswvW58
IJojsNdLQBsnXf3fQFgPCC40AdeZ1jCtOSzBnDBEb/GeDcgEezYSDbxHO0ENy+ltyUkVimp4Ui7Q
ChWivQz/EI/94O55maIVVblutx9wzTCGVXhx4tl7t2zsdm9ajjo3LXtrjFQDsFEJAWtzd33DIk61
tnRlAVVz65JuEWW++FDbjosLJks1IcB6+qTS53FCi7j3poZhG1NMeJViVTcPzeoBtyIfh+OBq1UJ
mttqa2ChWAS1m62YR4wL92SJXknC6wkyajxhBSgkTQotjDRUkF6GwKt0r6Uwm/FsU/VIrtNVU+S/
l1Ghvkm8rI96EcHYQH3YbYvtFP93uPYv29SlrFaaD8bfQ1nqynXhByKAFFpf9lKTCBHd7vtumwwQ
HqxfNQ+CVWIQu/CY0QcWezs6tkI/0zIecH/BiAGAO98vgkqSNDODSovcOwPLKSJsGbYOPpDGPC9d
XWlvQmVGRbqaRS4f1yiJfOkHfvSGw0K2a9xPqOomP58JO0qPx8zmcwe3zcWNuEUTo9HjDt+0vOuO
cswiTofx6OXehOeDkea6S6m7GAxCe1RLEo7iSBuf5lI+6GYk8MPfq341gfN7uSpxbNIOu76/8xON
nLCVtRW3DbWF7+7k9yv6SC8vpJ0hwulfkbNNL0DME/oepwu0VMx3mQEjpYgNCx1nujmNB4xaE7ej
HRGgY2Gh6Pg0SgD4JQA5evP5S7g6gRnwygfRmR5LJjK5YtQwvOljqcBy7cfTV59OOW32PRd0EQhx
mPGaR9kpjcAHgNFDmHOvfRiDrFFXOqo8vi6A6yw0PNWnnw6ZbCP/rfhCM7GrWBc9oG/cq44LFrzw
j7+XpPLWytpZi1D+2Ntim+PgczKbmqYvIMAXTprWBcZHCvOaZq7vX68On0SLLoH9bMjVOvVSFQ+T
fIQTT9l+iPM8Fz5CSB6uCopQMNgauvTF5imUOLpRyVUmFPEqMK+yl+GBUhEJ+V97wfdzXhT8rgKm
ywCPwa5VPK3U0zPRCroCU9iY8IgVsu2dD6nWXGz/lkonmQHP+zGseFRmCCJxLsqhesD06lDFvYb6
jQRpV+bCNUb6FI5+gFBfLTq81wa+CCpFLeGGJ3wiEecTSBoqHn1gXa8rH44K3HPGWoGmOKpyvv8A
W+vqDAUXQXvOcdUOyijW0zVoeGlPqpKrRZW75wYQmbpZK/r3v5Z9BPz+O2Jk/GaW8iMzMiXbEsXU
6hyI2M4dP+jloHhcSxk4w3a4dW3NeAhxhr+Pp3ejv6TUtXEi+NtHqlvlh2oxfODBNBi0pgJWO5ra
JmutZnHEd+Jp9PdfB+WH004o3OgU5fk4LJC30XyLRL+sVYSeO7oGMwbl5DhwOCYoap2Aa40RlIx3
mnkvhuy3n982MUx/CjOMC8SwwUxxoar8G3CBeCas3wLqtNXzIqB8P/IuRrZSV1cA0U4fQ7s9gN+S
SGGPXEyvBNNzVbneoQU3f4/1D5bU1RS8161wF851o9Ssf0Xo+FDl0Jofn8tSvdICY61RuwCwC0Nr
iKBRXa/yXGM8SV1m/+CUuyuzTieIq3HJzIzAH8iK+TH2u7ZDaGf7x9FxQpbYctsKcgxWLtA/UiAp
VNFlDF0kEzM/Q9EUv8U1Af8d+VbCVx1P6mHm/NBzec2ZDJTKKV6puyYkHn/xB5Fg9tWCE18pydg6
Si4tAozRoOiGgovP5R0qmjbedUMeZkaEJDy6PRZM09v++/Q/vR6hIuzVnj38hA/ur8xGSPsZvfda
//2DksbJtxRGvBxDJ7WLs+jbfCdFHLGx6aw30GNGH7YCYVlwM44ZVv0d022e/DFdwPiqKDyPCGj3
kCcvgzKTMcqKyR+jTshHXFoc27ewmzM3w0j0RnADDVHNQSJanPF3SoOjGUmcLrGfJBW63hHtla8q
PyRxQBjRrWyhFJqt1vS3kvwpa4Oxw//8XZbmy2uIEDCoslvKHn+WIgjJjm1HcfbGFT9tDluO6a/h
06fsmzI7F6iLGb0AobFgjWUl2fAIExGwRTSFaWvwLS0GhYTmW7KOXV2BuTGwPljE8ax4PRxz9tt8
wnQ3YjPoBt7d2mlpUWwHKqo3KQJmBzEDlYSO13WsuHK3Cs6P1s0xeU0So/7VK2s561Xba1kQFE5t
Yj7DKE9G/IAnL4omfR8zsu0/mfgtEmlRQpPzAcyZ3NUUXct+KUCDNtiWB7pQ0SBxTrLIGJVPTzEu
a/cDw5ezaWPb0L/YQNwcZFzXq9FN8+Sy4wZgsrZXZkaJq35k1SgSVVgD+HzbXNZxs/1Y9ZqfXH3I
yjmAI0AWDtLi61AbmiFIweUJ1P8mcKx79FJcCisu/riIw6xizNgHbUjyX3c9tDLzuEOh9Lb9MFun
wIU+CDxZHmMpIfPdKRMeisf6vqRFusqI5MQ8NJmF5Bh8zlD4ukY0o/qhJWztE6FSoCNZ+oHbqx0r
XXlQ/4kxQO6p98BSd/vfMSKHzc81ti3ki/fhh7xAh6XP045jpcwNBC8zU/zcW7WlaNK2mP6tHJpl
pxFybZSeTXfd9Ofo9GLUQ322wz8SfF9pyuA5ovSC+FKXnBojqYpPUC7o4hvp2oIk6VpVVbkpdzoy
ortTWSobCtj4+d6IQgZyxDcs6lWngtuxb6U3CNI74BbPF4EEPPWx3s42ZdBUFnAam0pYZbYpy2or
LewVn2b8Yzo7+zm3dOM8/HwaRm5afA04dFFZvISLd65JCEeMDWMs6nZuksl55ee1HVcrKvW3MqA1
VvfC3zK6q2RRiOcHiYp8Jk5fltMowaEM+MavDzR14g5FXzNV0yuC7ztKNLy56AvEL6Pw9Xh+QKeQ
xfN692H74yJLExkjgs6vpfMNWOJzv7fBMj/IWVEQZmztsOYYjL1CAahDY8DKHi19gpFXIlTgD6Om
vwLtKA14S82LweViheQlwyFzgMZdIrqr/GHOxEiJpiTzk5TbyDemcT5Vue/2zTWUqOsYbAo3wYeO
reZFg70/gLfrm58NkzG3aAeEGrAg8GlhtKIK/FgcDc8E3ge2DmGcBcjHLfqKM9i85mYzAEE1lPd1
2kCbgYw6dfnRtTRiaKpxFM2DHlFXG0ivrFen2tmJS4PQO6JCjX3oecqv0HHhhTzIow8kMgNAR3Nv
iRbSzIJOt9HvoanLwccmF0MjyKoiipOd6o6+5agrtACe+kgagM34MFScMQQtv+NEE5kKfFDEdZJz
urMjigwVP0ihLt+vQM90vbhImILFdXr7wFqmw+S6t78e3dJU6+bVBZNNwD+cHCl6jb90bU84GWU1
0oXDJ7gANORYdIMHSfMP7JrSHzXdybABIhd0GWBM2IVcrvgMn52pcihRzYGX0DQNk0DvK9PSLv7M
/bxg0dd4bA0B35PxwiIGb8DRO1Np6BeaYRJ/fJAX25jW1ZtOxxee5QtoMrIdOt1YKlxizqSqClBf
FGI17xZkP9sQLXZCd6LeoVGphnEatil2uLOG/8TtSFsDcVF3sMvFMNt3VXqY5u6tmIzPyefEuCoh
Wy+GkpUjYbZGfFcHh4IcBAa8iLHGQA/9zpg+qNL2sHOsYwxABxqlUAqZbfyELOB2ZzklOJ07sVS/
TEOQ26dLQ1u9SCwya7FkNLlNG6EEoRdJTMWW4eVIzYTx+lofKAZaXvc8r3QnFAJKVhXZzxcPEj0K
xS1ePLbpDOe8cGlXejSFrzDY/HhmVSPeNLPCAMWOpj4Ng7D7iYAfne+eTdn4WG9v4ZmUeEQIa9RK
OtfXcViSKCoqvfm+maTm/IxaBtZl/4MhXDGkYNT6NqeW2XK0jHjz11ISRFYeEZtHuWtk/sHIV05B
HApAjHHIp8uB7zdFrDXXUJLM7cSJ2krL1pqYJnqpo3inrGnGDRsxsyV9mVE5NCVltPoWB7fvIHox
nNHaEYnt53pViU5pc4voSasjyoWsCYmXTD8X+0HB3UXWBYMvT+e1y+bZPlPFplbdSeWPEa2VKZjp
QNbAtXrrvzJO/+jZOLyiiClUnUhrLRgtFl3g9sInGqy90Rh4BQCw/gvTsNIzcRvPcV/ULZYMoDVZ
Gm4dOxLLgTmo+Oy3KQPFmpcRTI62VE1lytIlBes7tH61+ugd2gUSMhOu/3MTKbRQ2YT5rs7V3Qv4
oZGsQrmvIweunl5guuAZZdEyqtTLQVe2xmaNB+5c4XXLMD3PL+aSd5d5V0JK4JkMh98Gzz2oTcAA
8Bg7RH1s3fnBkKuy10gwLfEvidwNiDvfkqDJCdriogPYU5E6gXFvk9YwFHd21sZK6P6Gwp/JPb5N
n3vBiiXYKBH/FOTJiRTXj7qOL17aR9OoUuCTl7k5Yhzxf+a2i8rKjg+HYKUbnDcyUP5F8xsa2XTP
NZG3TRAP12pGC2GflB/B9m3SK5dwgcbafIASKlxqvLEEVp8MtYbg4a2wKqTk/9pmcFw6Knohr9hn
AAWNigWJ78K4pC5ADsa52qv13W7F1W3xqzRpxgFHfPdpPQwYTZcM6FttnzDlt94+hJF4xnrgWbN2
rax5TmiphuRg+WquiYKt808/SkPM5asbze00mGNGWAkTnh6KiMULoGxgdl4lUwI6lEplcbMpjIaM
v+PP1HY2MAhytsRRbKSOGKqdx/8A0g61wiYZjWvyjTeULGhWvKMDpgwiiRh5/c+i7FP9teVCxkKx
oPUxJo7M09F/U6V23hFtSVTI87Zzp8c8HEcaAdVl58Pcp1llB+xEBAgUOr53vvWygZ6cHxMErtrE
kQjv2n+CbATZTSeXLx5g6+mCOM8nZ9hmKdC1O4VKDZPonrblzkunO+ydXbJuDOXUAl4f1x7G0MQn
AssPw2HTOY9GYm7PR6ahAiaKF/BW44lA2PInO0QwvF3WG4m6EbokXFxsq8tnvhJKcFkKXje57aI9
ZiVBvSUdcyVRBuZvfYKYz86rF5TOIzB6Apv16ZC8vk4Ph7/ssKG0H3tSRYFZ5pujE5QxbOvaiZgK
/oTQowpemPSx+SrSYzekKfigjW5GwL8YC73p0nTv9VnHg6XsGRiS/PcX+e4P5w2d1KP5p+p/OTKS
rODKuaQA1ur+9bIglxPqNlvdPjx4Yk6fj5cRs+FfKwB3lJgstgNJUUIDUublBxwE1yrdHukNO8Z8
xBcPdfuDcvNCdeOcDzrzQge1ErcqT1Rieeye2xUVjQcbiGjGMQfJe+7fscKCSiEQ6SjNYzO1Piw+
yxuwgkUxXCesXZ23jEGZGV+eYIEUFhZlMBs0wq73xR5AMZmQz1pPwoWb3JbkzV+A7ZzkV9+uPmrJ
3mb9qBr+ezwdRH7Pbs1Rb+ySoCsaFbUlUTb+i00//RnF4KsrNuC1ZCQdpiMbcybbw8sTKRiYkcrD
SsFNctY0+UydCLdkFLe//Q6ZOMa/2vAC3CN68PXxlbFYXhyAqf1nc9z7PzkFXrp+i2BXjIVNAySh
ODVQZCEBEAdhZcMAjsukK7RkAfD2ZKHKwNX/YWgMk+7pGElkBPmWEeaj9C0ZepVpHExVHRGMJjBV
Nd45XSo+S2ROi1a//Ljbbp9TBmL6BvCf3COOIdR5weLybjstFE38aVq4EGO1gsPaS82NoJ9v+Txg
s9h3Uz7EvVKf5BKVm2nUviSdDvFDdv1xxfF/ilY94OSyb95I7xkmQOgefqp3u6Xxgbgsd2BIRBYi
aX3dJxxiYRQ4Mr+XLP/l/d6ENNr6TfkbKn2Yus8n4uhR9/FFiKCoFe4F2vFFnsuSlXZpDa0YVezU
tPvC+eKTQdbK4U9Rl3hN6YzZ1UlJudOeWrclDGcSVjYfnHrSCkowFFCg+IvqeoyicEFYqxA3Jyyw
7HH45GT0RTzF3Q0GmVHBV33NeMJDBw/OOKkEjvXT+SU+/86+PZ+Afg6UXcrjGrJ3yEQLsjtZaZB6
0xcuZVOthUUiYodRdud9EBIJgwi8vhXO1rIu3foyz/C/GXSkUBA8IVkNhzQRghklps/vonFfRXJE
jyYcn6ZGv/RVWTOYPH/K6C2bCq987YKK3oBAnO1c/dGp9X+Oko153oH9KACMToEYfa0SS4b70iCn
Wd//nikw/vySdtH8AIYj5MfSew46ZToi38MMAJ4cjT/f+3QMEiCRyL8fPa0ujDZ1WjwS0ORkXNx1
YnaRdb+jymNDENdMesSwR6Q0M5pP5LhI/YFJb4nEIRhkLoYr3tKAaqvHrxRyKqJin55FU9N+3D9O
tXbNmtF2/kpNaWJ5Bntm8Czwf6A8dmc2iA3e4TLuSG6evfrP0G4HN7c7hL9MRB19OVWSCS5RY4k1
PkAvq8cVX+K2dNn1v8XbLoI2uLZpleEPXpEqWhdMnUnG7TuDxi2Ge76RacjEmsAtMDz5YHTTbtW1
9GcD0cVRriHfmVORz5RRysGUGxgNMcbEu7sp3na7r+5gSEC5vsHwcjBZRx0MH4OLVlA5c73/Qw19
iAeBKWQrGULI7Bo5IXFG1YyeRlk1wEBio5PI005vX1WSkGP9/XJh9bfbAtmbPyvLQaHJxeCHfQ0t
ARIUf+MNXORkexFXJomZXN5JY8Kc1sNOqo1qAErKm4ZqOmbeFhERp+tphvmcJVzWirb+rZSbceIT
TSa1Xy1D84XTF4HlEWQ7alAru38oB3nshBCgIWxC1kZLlNAsakWrepzRRVNtfnEv0yO3oosIeSCh
NTUyB8DVH3DsTWq6yeeBeVaRVMgaB7SVv0mtDn3dIwyRn7dDJUoj5fqFfEEYeR1RsoNjjAoozpsA
64ERHjBMqazI8B2RMMaaUd3THPewXJ7zZmtHlFvjuSkSGPSbFJklkz+xFzh776KV4l3YOmeHTOLX
KvAJSVOchEk2io6goHk1dpbEERo40es90i2QIbe+lmQEyrR51kYYf5vG8UKD177jilCh4zieVywi
kZZtJ6iOFSxF2qe2U9txeZKSp+7p64kaUw3Ja5isuac0PmTfvryHyikTb0Yv8a+wOBfX7XB/KyIW
5uezOXCjSnsu9EtWMSt0NjF673Aj4NzBHtd0ioG5HUxWBSFbN8DiaRHS4SxnGNASkrSiLicuvfNd
ZFf2Y0d33sOimODkgaWgQNLM4Ax7KwmOBEV/oKXG5fS+xMVCsip6ZsDaYwa9SQjub6dbA2KeoeEi
Zecd5h9Wk7J94LM1Qbn5XiqsNB4dfTbcSsLJA28ejDuhOxH8VDxAB02/HSMZFCBJ2CGgCXT1tTkU
KIP7dOCn1tErRPUqsfFyvBhOivRoWy0Gq4k2zdiUCVa9b6Cxu9VRfXwNqDe1YiMKAyIQMTKspekO
xMCltF8QV4/iloiWaKP9d+CcnpslpUSLREXUaNb6wUG1Nhpw2AOA1BsVLM6XT9++7vijEel9lvRz
WCBOYW2ZZYK1zgcq1Jh3bwqQ3BeK+khpiXYLUQAXJ4nfjh0jL8an5J4K6w2JUmuXs8eFhOjPuIOf
ljUEWd1JsoLtufL2rje+AHQ3bwDLvv8i3nv94GGKkPrsV5dLjrGsrh92HY5Y+rp8/IA0sFOLf2sb
zRnP7NWUgqfNzhejTCQGVxiF6IWVJASK+ovmaRNiBSb3qFLro5UhdbX3PmUqFVtfhLhyd7soBhA9
PXNXRf84JaAB949IXZJkUn19lG/b4vvIrTpJHS4qRsUT5Kj/cFSEu1HPjDWyXb6MJlM7vKDi9KRE
wsAYWy7gEotNPjkvEVLUWfPcINNzqb/c3RrueQ7e5BQIN/l/WDDkt9r0Uykt9CAIkmeXRmtpUSba
XJZQX7sbZzmWqoxtJmOSOGyZmPIOUxGTYTTQH53q0gjbA+JmOBDrQFF/HCisOIMfPss/w5HEjihN
Ca4h7Rch5Ee7m9stcw17wLEKATGLwmuCROq78bzcuOzq1pZ3Bbtu3iZxZ/WWmlqydsq1F+rLWswL
CSa8SvX2lTep6xyw7l8SIrkvUdpIBCZMK4r9btq9ky/m2icf51NcQmtsCGBMvqrDZ1LSrljWPMC6
i4iH1YHlwyqkF3uc8BX1wRSl13m6gyYmR72whuUky9CLnRp5kq4tnAitUNNspM19eMzmAPZFDKUi
Af3wB2FZMEf6nRXIhhUhUeypTiyHsTrp85Btf4Q5LOaJahgnmH2BRtz0Eef80zvoUCLBrZcjsv38
ByiKXvEmV2Em+eWxgaGGt3WB/Jb1l1SNrx3CIZNopOORSAP9fWaGW8tD0NkoVSsXSXWdt4oWnx3r
NhQ/0HmZCuAoYqDLXfRsyjrUtD9Kh3DWRrgWzjmplmEfi6wbQBIHtikIpVULnjvUNpv1O7hVO/TN
+17Jq+JG0RZ8bjfrsyPAlnnO7xQOJ9O2O+WLXyk2q+QfmH7/q65gaWvjk4nf/sCQreSA8umBJaa7
nspHE50rdKe3jLwn8aq+aXXOB7ymraC6Ka24+hVULs0/uWDA0Yrh2MwgKTH8tE8LJFJvIhU/bPkP
RceJol/b+1wTZYKBoExNcVtEeY3KrFz6FZluXNPGqvB/Mwy0pqwAYzfRdTRnovJvQutZ5cC+XoqI
nGUBls1KSFq8vUwyRiJ/V2jFbCC8M/rA/O3hiHjM+SN/cvJb4cMO1vjMCUfwa0VEvmxOxF4ehWpG
FvkJybgeokwiDtBQodVsi0mkibvpg7l6LudWPj1WxHvESi3c/4VRJlDL8rdNc46O1IJEgJhdpLFq
2yrccsB0qsYEdEIlaupD1wtEwSsewgIsjT99slNYDo6pzTW4MfOT0AmQog2NTQ9GkGrFolP0ysrd
MbRElwiF8cJvtNfR5ELFSIRjuqMrqwb9i+EEDNKhalUY1xU94TI40iFZqWCUhy+m9hEBWhWEu7OX
BDL8/W3b3s5Z0jSG18MAJC2e9xdY9vhisi5sKWl4no0GT/NthbxXISa0oJbQ7ntveTz68XY3CslV
yIHgNDqjZgj1f+nLAIDcd6VxfdBbC2eg4p7sa8uzlAwKv6gCF97nMQWweSvkaiMWUwmEPeSwi2WS
Hp6nov5gxArg3lymz7jIQU5i+BCOipdOpjnuUqk+bxm5sE/Cl89bi+fstkpsQ2r2hVLV9quAQAr9
cgq1jtOUHUH7qS8sqWD5ZVaWdLjAsPW4JzmWBZkVQOgK8ku2sQ86BFKMQlrGYUyeg1Mybz7XTzvq
yrMUxheJN2e6ACafgQlLIj0t1qPhotUsW2Wh5GLylQFAT6dfUfBQuERe3gSaD76vutKnjaNL6ICY
wyvEu5DITduvobAIoz80l3OzGa66rbhHDaa5/LOBM00RICZYCOq4Hxpk8ZIaUULemKpMQjaYGjwO
md0/kZl81KmNDRi0JV+F0hsA4c8dfDMr1FvBeaAchPX6MRy+eBCTPItpjNohNVR+/c66I3mBkdQw
eY7M93bLkrDcnK+EvE91uHcX8xs+wBwmtOrozcFbaaCvqyCMe44pCzXap1COUFNAutTUHxbB/wwT
yJuUqZhzhJw7NDarJpTTHFSEm9wtZ1ftj+0aYYxHPxYUDt6SqUT6VxY2FKmqiczVpqdDwy9o/LQ5
NHiW/xI8M3aFmRxk8ctnl/9XTlZgmQh3pgDeMh6idDy+axtKb3O0eerfrBnHIdnnnQMPQTAwl4KL
6cXLOalZxma0Pv6VEoZmLtpbVmc3fQUIRiaBlKTRINLtKySbfcjfcusGBR0nzHoJkL7iOBGiIcjc
lsWU/8pw1SWEAKebLHu32Mloaf+u6vuOTTDIZQJpUPvoz2e5tnpCAhobvr7JGoSYvtup5/bhpQEt
88WHp9+FO/lLeReRSV+slvxkZdaVt5Zyx7rmELd2PaHkhxGFVmdXV3Lu91yL7HBcwAxKFVUK//cR
PSjzGgdj7XqNqm28IJFy1BKfbwRLKWn+bVTrxy0nFWuVwDKONasNeI6GRdeBD9fVH77zAMkMtxbn
H3o+88OyKMUg+E574cWX809I0+RBHvAvubD+D/XdOdGIlE9VanzW8f61E0ohFtvnc1pPbwMbuPHx
ACnuGu7m+zp4pczB5EO1KjJ+VT+SMFhIhZJnQdnlvwV+46uR/2Dc6DKEHtGzLs7BUkruEts/MmPJ
MnOsBA2/au03MN5to6bfi0K6rbF7WkuFW/GEDOrxKG+8YX+VQbPpiMV5yCadvrMrRD3ER7YlQ+tD
E4PGABiyDqcB9R77vthHP8+OlqqSlBaVUbgO1ZDmySLqEG2DX1uRVys4VKn1+4R9BdR9FWkdPKwh
Q3lwSUEQtxHeNBYMi7nNjyxHK8GOwdBVTNtDeorGJ0A7jzW4kcDgYRACxTwN5+qgGfpADovhXoP1
AG2WJLUcnDlzXa3diaMlF3llZywEjlf7PSRb5pgRnkee9rLPrfmGd07th3VfdaonEManDJx7fusB
bsPVypZKhXWi7FIS2LKQl8Z+b6w7X+ylGsjD9WVKKaZGlxnDAGjvp9iOv5/tdSyscjrzb71wxcll
QwDUoExKfZo54wYFKfHTpNlKRY2khekTFb35QTNUCD+we1IsEllJJ9QswIs18NzVEDXXwjMWYYTW
Zjk9fYPdNH+CE6rea/ZLRVbkbTJ3f9/q1cNOvgNK2oXM0qG2go4EMkbpy/jemIaZiQv4SJGXTi4y
ilqM5eLD+9Zve1EvXgKg8cOpGtE6YDe2OccNLBbBT+gxnRGEDcmmzsVmWhjZ6UJhFF8gWqpX9GRi
71yn6f9RfH0tZ0qYgiJayORoBjSLaxxtovpCWW30mN0EBvME0UggxiU1YyElsaWqUCUVbAZ3ZOZg
ceMto1yamxV2x4jZ2oPUJO6oOkmJJTAGigZpEOUlMgb6h7DQJyDA/+P17dUbqaP6nAI21MSFA743
mWO4oPDci7T3SP3v9l2k+70DsD8fx0UQBZrLeBRRdNIHGBGAW6GjyRb/9LNeSNbRQLNwwQSSa/ml
mJrfcc8INi+1plwhGxnI9FWy55L/oQ9mOce0ASAGtVd3nNQwD+pm1bYyDE5eHWNmRFXbDm11SOxv
JGptAVK4HJeK/+IC2IfqIwg9ZZJV/yFii76oDvnrhvvKcZqsSb7Ef0DfS/MGEf4DBBBi7j0HN1cf
0oUGwzh9MSPsx07UDxGU7NM5RpSsuXcTNypmMRzkO7d5zrCq+RniH0vHu8mm78Uq1ajVkj91uzhJ
2DUjlNN4t4dTTXZXdAEKa6z3E7HcySxcRrvXfopOf7rR7V1RQAZyKJADGqyhif7vKlPOEOn83f5d
OkdQouU/GlFB/4nFsdWcHpYk7L3FLgmzTYqtMPCH6RnJIfwEM9/wOCY5PLHsyKCw93oO+Rpr4Zeh
gY6JOeO+eI7dMU81R8Ok0spZKvoTHFBHq/ptWiFW5ivVxYwXSm0EBIlx9GzfYGQEdJLNgnRkzHeB
hGNF7Wxik84y1UKbpkdjDyIAwhGWs05tx3TZcgrTnT2BWaJ81uc9C8n1C8mCs7ozXSYPEoXnfq5W
/Lr3xCsux0vz1VdTbzdpBlvoS005j9yWIDrkFSEKoZ6R5LaPVtJolhDGV34qjHHgAl4RWPBltl+8
CbK0bL//lgQFl5iy54LrfPckijTGdzBepPiMK28q03oXinuxbAOq8PUG6kaM7kqiyVBieEts/AZW
GnPti7uXL+SScbmRbFSkpcfafj8B+0YJ0hECyOvJkCTGYfOsJhsqJjzV4dbMkeYnLRuK/QEthyCB
hSKiTSSnICnTXElr/BbyiXlSBAIMgn9ctFVBoFp+5w4WLxslunXf64spMfA2T3H6d88oOo+Xe0cK
qaxcjCijYkVgVQYoo/h7K4cjK0phSAVaTFrvwi15bsYIY+TWH1A8J61jD0cg0ERqjYiXiVUP3Lzj
l7je5VYkjuYtT6MXVY54RYYCxUFdAYQDEyXHVR1a7AEspHs0ZkLSXItyNxZCBIkVQj+fFh2zjTRE
EXK9HTvPaKd9wDK7Aw1H1cDiRcNsNTFgm94Ihh0HWWpnfvdgcjyF7f7RpTc0cWG3gsxWApfr9dfD
9gqts74QV1Tylxj6lI8Ke02CQaz2MIc6kqJv4TS3AVkmFAG1KI/00BOp1EOEQ2hy5+hcIfXiETYv
TclOSjroaTRYNjvXpDD6PpHVXv5bLJ+hk24GwmW7SHN+YkHeKqOj9tLIB2DGfZ3ewSZi2ZUXFXum
LtATuhRy+JSh0JiMYUMWDJU+Obf7ZKaib0OStYfoLkxZmvVZbjPX8Cd6VKk+8tI271XyztzCilnl
BuRJq3VTvFBgBCrZO+AWwtUblMxELMNs/zPXv05IiyrmZbu392pK/TOMzUCUOagKLLSgm30vIrI+
MnamGWhBuTgQlSBxFuGakb4QbuO5sTqN8JGadOrUMSAVIds6anvsrb3wfNBReaFJCrUssej8szZ4
ldI4TOYkf0QoVuPKim1/k1O6NtJRFG68iitxiMC+X+30z4F+dVv45RHm5VUAkX5JG+2p6XEK4+Ug
gnVSBw9aWUC+IF5+miPQl65eIM3p1fEQ/TM+0Euk8BW3Zv3Sr9vx58g8ypuVhj7l3I/vppyk+Ts5
PDeyMWEH6Iq+CrXxhTy+6MllR6CBt2qUjS0QrnX0YwS5a44dZpqGBdwffyR32FE+FlqN9mTFcVi/
xw9vt4lrkpVgiaCuUXA2tcmB+a2EUlMBpysQ1MRDIDw1+xQ1JGcggu7Y9RkEMv+iUaJuyUzCrrN5
WH8JFtHJD2In90MP5AZr6qEC/HuBgK7KOmj60nbcf1RnqJErKmVhDapa5EAL6ZHh4a8RuPIhdkze
Ttq43TqVYL9i/C3wZeV2+DjtPqgpQH1aG6lDHAhFHrG9s1oQS+e6OP4nVynoiqimA0EK1DPfIr7z
WhniBW8ib0YBPMX6dHH5mD+YsG0sXc+Lc5kC6in6GdQiNscvmf53icGAHRC4mgePwfw/O5CEh9Ye
DkFucO/cWaJpb5u71eKbQOP4eJlGV+rQByl+QepQg6jnWJlu/wUwDADU+xV6o9ZXC6lcuHO+i0sh
A3HtMrpL+m+dQ/vmqTzd1aSei75eCWCLeAUkRRIwxNJvkWTZuc+N+FHl8l1vWyOwvYo9ni20HzxY
mvZzDmgH1axkSyC2urJjsH5d90Nodh2KOMsELyP2vSiCZnwARMPDaPhlhxRZUXpSwXJKte6y8+QV
UuGTprd8kexeUpN9iA2UZYMMM2Py9Ypiu7OwO6PFaLXl3evoRpXeV6wnTrEYGX7Ri9JSoX6jqIfK
h1A9baTKKJjXBYdzygG8zWlMP18FBsj1ZVxU6ew927pCtmi/eT1+XquEFisRocgvW+PP6bO+t9cg
1168L+zpkf5BfFWK2a58ZP77RGyvgG+8n29reORMqxscniawoOA88gjjIeCnhChEg75jFpy/wQCk
Hs+OqrfVqtr0OxDY7nCJn0Kop3QA8kKC3F4hIPZxVofISfjdEnfpcPEEJf5JhhXPuUyOatG+DZ0Y
aEY+MT/oneYtL63zsxMSUVl/weu2OZ7Ca9USmOUx4Bq2DvTrQbn2JuhZrssy3E4U948sgFQPnVGV
tSeqJUoW4tjUFALrhmBSCDdktbdZsejYh9sgorvF2Yol2x+eWqbvWn9sxz9bToRadIFi0BwvZG+3
60M7hjQ8xanVAkWiUidkY/gZD5u+wPK/tGzvZxkWkr/Vcap5xOlgA8pB6lMwCjHHxfO/OSV/tjVV
bCGP30Sw1M3kfq1LvcSaTmg/63j5rFZNsr+Woni3dExhcVx+O4Huq/o74c3mnUoA6+nWT2i4M4fL
rii9u2Mxk2OgRZkYLogT9N6MNM8gg6VRPW3l+GPuM5idzRzXVnI/kDNeW+gUMke/4G18vEec2CYD
X4ZeZchgnVAZUfgaXVf8KLxTOAqKFGKnf8cza3hWUd+4DGXBVu2XL6pqeWxpQUOseiYqm4EVfpjm
48j4dKe8Va8QCVwn2kPqxXT4X27RjB06taBkFyUBQglPuvlA9gs0lcUCtNe4Chg6rllv0aLMQV+P
zVCtO7rT5G2vpg/QU3kw6TQ0Nsk+TXXOunCxkvSQXTUwEJdJhWpVE/NUe3EUffUHXBOci0f23BKA
M81ObmvVXjvM0IapDOAk6lzxf9EE80rVn1x2MCsYVjF/kQHDWCKR1i4w4c9nVJlUEgLvxm11ewUI
I5xXsNp+eVWfjSIn3JtuNzpAXYNy/3jD1NbR+c6WE64G5zRnDXlvkq14YFDh4BxhutvHzWoeFaHV
Mkdk/YUmeY9FPJLhuFQMNj6dIfVNqDd9XkPhhng2QoinVWuC21qBHVNzaBaB8pdTrPxcltUB7Kul
gDpvYo5kiyJWt6R20KPOIEux/lwtZu2rwzyF1Lp86a3dI1W203bDHKc3QxD0r/VM0Hja9PAz4JNO
IKmsBfGbZDTOUD3t9dREwDFXKOIjgXoMukztL4u6RASpc1pNwaDPAP8yj3tWM0jREEnxAu9s1nWc
0eALYaIwGjApImkzQwU00ZAhDuMx+fSvv5hiUzBxd0fQf+C34hcNziesfgj7a1rjqTAmr6qc6GMH
ZDOE5u90GVE3qCYlbfh3v3rvwBFPxLpyvLy9uMZc15DW/A1Dos4GppWAdWOVvWqmJ44W+v1+4yXX
z8iXe6m4beU8mdT25ssRRfj0M2KUafSF/jqxlwCSybR+OB2DniwXouVGmSZEo6IHZQ8zBgSHdikl
IiqCjj4viED6D148fbkJyA6eD6P8xUg0NB0x9zL/anadY27dYXyHnghwVWIpnrTYgZ9aNIqsXaiq
OC2/j58HVL5Jbw9eTBVsqE2jhpMwhm1YO/VnvfVWCrnTyyBZ+g8Qi0f0avoArHPt7Y5BY76oCRvz
A9oTaVSh3Hls1TPwKsytAMbbsdD2Exy7/cvdMS94EtvmiJyvoqbhA4yhyu4xHXBVlfTDvIyz7D9P
UkmnhuojlxNMiQm5jZKU+MoAk7l5TxvR45SSEQs8bCqtGTIpPmeSsbC5JnVqrWBOZJaID+1ReEeP
BenvpN0aXc1eB0Qijb0Ui7KbACwUkVHDv7NesbIE0nZdSe3Z7d1dvGslZVh/9MohmPW3kZe/C5Gd
3o9+/69P7GLQsUgGsZffux5RkQPqUAuWUA1ZdE887TA9ObPDbJlKu2Z+oI+QXSFigidkj7hOWagV
cj/AGvVPEZCaUJqPrQ3LVtUcTsrykFNvfKN+UrhOgZ7HFkiy3F5lJ1jih9NZqjpCsmWFOkDuEXRq
jR7ZH8QIZeOyDjl3700uMwoWC//umxWvLg4Qoi24JJOZlo/hbIPKUOhO4jsgkgu+Q899YOjXQWfU
QOfpIiEo+Nz/Lrbhak74wdzEccZ3pxSh9+t19aCgVqtxsaoYFFAH618JZUyoRSiJcf3c1sLYOOAL
iwRLkmxhjqxf9i7HUZs/A0/oUC+C5nRDOTMtLFnC6fw8RP6wBFh5p5GNBPGp11QvtiAbnPoLvfCf
yg0YNXJKWTsN/s7x4MqkhzSO1dlAHV2fIQrcbNmMm3p9HOoalzAKcWajmJTwzNE4rAAjAKDJrHKA
ZNjIrrCattWpcZIKqrVUyQ/xoCwVw7e2QYsBMdtAzflF3385oZgnbM6M3TXigKKnNx26sOBSwbNW
mbDgA0j/Q7GpPnywra0OFsGfzVZoTPyigCOD/pLqFvD4r+dnK1ThtnFf/oM6CNl6r8+BrtmvByfR
8JHmYR+IEj8VFHuF+nMGKt0e9ET3kd634gRFBksgx/Jc/5sthNG9xYHvzanvtuDZdvDJVP+4L/qz
GcLLh7hO6Bt4X8qjCu/5TkUaezJjFQRcwjsSLZtxY6wqQcHDiavdn6+W96F2Vd41QJUkpCYUIbMg
5TA7xIQsHtnzcdf1D8Y3bUCiMrpJ+I0X/PmSZ5Jen1SfmQJn/MyVyYZPexckNeV/rTLov3iW0pXI
LaHxMxUkd4yhSgIT6CVC6ej1bSpgS73z80KVwi2ERARGDRvK7yi9xGI2rSp/X/eUSP2QMD0KmKzQ
rWOtS6wGPW80Gb5WIBaUcsjBaZCbAD2wN+JnWJLXJHarYZuZpj0t3YUPMOZRhJWx0fGDbZ07CPw4
oIJgwnRnpttGWjCVDv2l/5jFiKPx/7QWwTLJCkHEt/o4jLRSCLr8gU4kRj3Gt5ippg2Oc0LHCfH4
iJsjOCagYR/1ffxrqB/lmDnauauK8C0+/XeZgtiC2CKssBFUSl+NcJ6pqZZLlyLYTMD1cgE9JACz
Igx4BDSXN0beP9l+m5MY330MN3DzX756KyVdtCVrb3H7SHd8rcUe4rCbQtbfaF3vl7ozc+oyoCU9
AWrO8azScSyvOGPuQagtgj73k09WW5QDboJmZ9S9+mFlzQ/XTS/IAJDP4/n043tK6hONn2tu+vD+
q9Aq/sxQXIubFnOh7UEsWulM8n8R+adrzF9Sx9S6pyBfpyebp3Sh1g6DuokTJrZKVhp3qgd14GkF
SBSNoO3YhMBcdhRVvMicYu0RU3D/sOtYLfTMUOgK+JJy0PIZ2OIye6gNxIQdQHjaJ9cmduoYrVy/
W30zSIUm5jgi6jKMYLpZ8XLLZ/n7+sm+328rl7Q8+wUkOwC5OyoW3KBm5uynr1mmP9ihnFPYnQM9
TR7cgWN9ZEyw0qz3t7RULoZxQAxeKrNja9WzwjyCzR2LSWFaMCpO/Czd6DPqkSIuRWAR+A1YC7Iu
xxbasLs3LGCatIdLvMgTSYcQB+hRMQDAcEFvVsD3W+tk4IIv9yyur4ejO1lZXfRbp5t2YyPX5oiu
JP1gmYYah5bYs4pASXNt4PxefNFZLYSVMX77jiomepPAc4vgV+FfSFCrej02m9fAcwb4C2kA/Wyy
+B+h3ql0BWlkIL+Am/WVhqxnS9tq4/FJaFzRj995YjWZDbE6Qgy1RC88S1LTMac2OTRMWXQr8a/h
u7mJY6J72hbPDsAlLt7TIPXWRQD+c9edor8DZCY71ipy1Z802IXn/SERlrT3aJgDHQFXLlwwNcMP
JKTeY+mgW46L6KYgeNUStD/Kkm4VPdz0hphuqWet5LPGh0BcPIFNICarFZH4U1GzVHDQPPaoxp/Z
54/DXneYR6MhTC3/V1yP3plM218te7WGwwfYcfuIsaf+TP4XzrHC8fzKjHL+0nI9KXWsgMMPu9ck
G/e1se+TCiIJhbF2yFmp1lwWufftnkR5RvLf33SUyhSaOsGWT7FCySlBqWf4B0xtSL44SCacGbaT
2MXekvmqb138uC0CMSo6GFDkpBbbY6xH6jLFwmMTmEdJ4eooFTGULa+6c3VMaBKMq6PFoyKd0gMN
x90IUs7wHFL0Kb3OFzGv/MUbcOE4U1qYhr3LKYVqVzPUAvRke1GMnulIvzqqxvfaXuR9NP6v0Lbl
r9Gy05t4mn0U/pYANKjEwyOhHGQVPRmxhTEalZp7C/uxxaJd1WIZNbGSofwsyWUW9yUmx03kVr0f
kKIsqIGmPbd1LT4Z1d/hUT4vZXkQLVw8Cmy5z+NioatDvUTVkz3PT9mhEQJi80BObufsLRPeIi9M
tnuYItaX4YbrdyZd5R3MgOJ/crj2lEGbTPwyBkQxmwii85qmUipGYbFWzoFE5M/tmC2atUTGfZwV
kJ0iU9EtMp7cq4mn5mB9BMK4mZ01eK/QZuVa4ipuhBbxvgdHVV/Xm6Q/Hm+kN3uNLjF+GgIWME/i
wWmBPUoBBjbEbVKuZ/xNTBgDorxNNuco4zAboHoK+FdlWljs0TWNjOk6O3ozuP2U1iNq3HOMI1RM
YMXp3FTquAQK43BVe6ijCx9hGtDqkPB5LuTjwMj0AytGvruSpnz2Cn62Q/PhD+EOSsN2E45RafAH
SdBUkZERK73jDJFg4bbEeH7v5FRgDUj6wJh6lB7BnJR+dpVxUIyGYA5h01bjIQ7Ck8Qmk5j+EudG
sEhCQgZKGXmKFCXgUgo0yBRp0pBPkXCGQTRhbvpnmEM2O2iGuNqW2jiWuJoCqiVP+oLBoCMCWDGb
US8gKpK6nESSKcQxkwtC3mulGrQOhYU6B/6MwRP+UyzAGLtuB8nGMV6QyEi/oiCY+gIfdAz1TZ7k
4ILtNNNVd4xcBW9bbdhgeWHxBsUlj2E4Q7lveJiFExjUhDfbfljoyf2vmk50OsNADMeAU+KEaKpN
Ja1UL3HShMKBIc/iIxMDERIOMKdvyswKbH6DFLsTu/hjaBEqWlRfMVLJwMMjFMatU/F62IR79Y6C
amqu+qxjlPac3jJJ0ZqfGyNwX1YmQarNbGexS0aB+sWmT6eJdHv6veRy8pYXS7rH1ZFbG94EZtal
YM/blynGwoQG6aGFYgm+VWicb1mi9o73RVvBa0/ReAAfRGZq0w/gKllf3fcqAglYiMVdSuQ/OkIX
uzr3GMT5MnGCLtaoTQqgs5ndsT1G99JvETY6WaexsSJEeOOmEw4f1RTzOiV8FOgyUFdnf6uGI2Q1
s3FE/n5uMtlzHYc1qT9GZzxISv/P2dlVbK3ea5P0zB+g9WDVexT6i0trxqNTugB2g8fBPlvF5wfZ
PEcGbONpoYlqiuY9WoBwIxHOMl6cwptn6Cd7fWuUeJf6tdod/AR05MplmQEfx6TFByZDgglGC5ZR
FeB/xb3cerHzSIFEB0Lv30A+K5U3hU7T7H8kQkubNbXmk7sh5tuAMky7hzz/ubVlPTwHD8L8Pljn
oiaWLQk/txmy4adP0Z+DaEw2+S3GsVe/Xqueb2ArZNoM+Ucu7uJsw9j3QthMFU6Q1pzoLrxc6Q80
Z2iU4Y7V4qpWjAtpUIowaYD4rMRT9t9VYVUm4+sAUxp4cnhpNEBXj9ep0hT5N9f/QMfFTl2Ecp3a
+MdMUzPIl6wO7cDY49g2AiZXyTq+qQ1D16/k7qgHPq4sShcsxJ6APPwBADeMazIHu3cy/72Fj8ZX
wGlognwxnZH9SJzG1fu7xQdd9oAjFdWvMmg0il/j2flXkJWhbD+CGK1FwpIUwniW2b+byc5tCMcr
M8LThBIIfIZqCmcZIaanGl2QQe/UKsaIig/9we5kt63cTgEgYyDMnqHcPTLiblhY38N5Zch0z5aS
W29OBKUvJ576vmAVQTPbaPc52de4H7YIcRoLurnldWgelYYZHS1KW+s7TIv45cr1RIx4nMBQEbn4
ViUsrEukWgLpU43pALQOx4Q3uM9l4t10HQB5Qr1iRKzoH/AaH8ExpQ8eYgbXkD0GxoBL/DV7zF2j
5dJWyjhNr6tBiDZrY3QX+OTf0R+6Ti9iwEFqGDx1kODoCFVtG1k2HefhMjOoauCIyXcv7a8E9Iaf
/0HUHE58yhHjo2T1XRIdpgwwo/8mmoZ+aOGWkJwZzpovqOofNDwXtaXQ5RVlRtyzcXrEkicf1uYQ
OMyU0cuH/J/zfcWVVHNDmMIGj3Bm2Uzx2uyoC4ML8kJIe7K4NxrJ+g1ykENF6H+6SJ9VnJwWyyWK
vy5z9ruwefVMyWOyUJKXVD5/ittdI/DkNeleJdwmAhunxkS3v5NP17mnkR4dBgRUUYmQkPS9dr6j
bp/Zrxa5X58PxGp8IG/g9Ujt2Whf83gJ9pRbqz1ZIfdnx/3e7Uq8WyfBpp9++qpWr8qTr5+4uokF
QVzeRtV5TdNBCYS253SiUcoAAjuGlfpz/UQ9zZWnsFdQSBVo1ky5noQevE4ORhoQ9P9EraocR9vk
iMDX7W151tY1yyr0eIQeTTfyUdnaVmY5eiJrRl3B482ia0mUR4VV9DRAsKAxi+sABXWR/2NNQLs4
IyPdDPZZbLJkMp3FV28PG3VK8+uB7PF4U0ITxtVjcgG0X6Q1UHUagFlUfCIa2kWOc0M1DkWw5EZ4
6XtzQt6NrlVuye97Qw6GyWd2XhCa9ZI9mZAK2b07csMd6+F8lB89513pQp2LpKeE/SqPv4nrF8PE
5k0OsSS+bJ4o5UmOWVWsik3bS0W4FhN+BB35SUNRwaqwzy/QSsmP2zTjiuBFZK9LN8DJxM7mw2LS
IQeJxxM5A5AA78PNXN8svkVhrJ9rmc8ic/IS8uZ5Qw83Nn2TutdgFqyorhhr6nBfYz5W37DIY8E0
pR09qO4g44hJ5vzTkDXASCkUQakGUyaLHn2vVjIGl/rK9OP4OXSAi1OFbi/nAaomts7IY6rY5xMy
3haIBe9THjreWxxxHh2pkas0xRxriXXv6usHZOzAVJ5sV6lMZ227mAXC4ljA7a/wvs2wbqeZYo7w
3xo92+bfTvWoNFLTg6oT+CLbEYyGl8I2V0e0qXaM2211mnGhfRuoasfWfjrrO41czX59rHlSx4wX
75qrIOfNV+EQfvs1Zyn8c10Bqwq3mDbTQ/HI+N3ck7PDozZxPLYRiGhtg12G8QXAqjtZMP731Jpw
lU6WkvOb0uE44gGiPNj8C9cZnlSszPGYkZpFTyDBGF3e+6NIhzFWx/FfccXfWOh+3OvGjj50ZEMb
7YwaHLbxlzzflecFA58jsYde5nZMLB2ZGhjFL7ckP/abh/dtM/1ArOIQwJT9Drbe5biNtQapBeQQ
3IBlLtE0cwIvXgO1r9ndUEc+2M7CCRM4yo3FPK9BQhi+b7/vO/Sn/u61lJxOl3+l5LNFbyiEWEKu
5e51p3ZfOoKAx7CeF2Gk60cI15IDxCy6k8BEIh4Q9erOYGEdtEsqRBSpNUVB3MNJD32WDKURqGop
bcm2tHetrNsdH1PT+79zVU23WEPi2zGNJ6VXP20sfXOjpON/l1RJLCfPBKIXE/r//CsBYMa0Z1RH
2mFTiu1Z+1d40GWMGgqGjUwy5kmVIZqeRXtqswqmnWKnH58VUDAhwFUM5WwGOW0rrN3PjEAgZCkM
myBHF1dWLOOW5PFN6xQ7XJYrmxUJZCazjce4yfeXxBQe/qffb+GgjFnx32ycWAF7FA9ORSe/MUMP
EIS6LhgGl3qzygvfO1jH2AqjA137lO7cafop8xVKT2bZ/ttwlGRfuPdO1A5CXq5SzpQGQedOFpn6
gKwtTKEvZsuZeFz7FTJ9de2q0eB66K5si0X5xyhJfJqqcif5BKB4EqxR3/EHxLWWzaMFPOuVbp3e
hl+aBITeZADI6Wk79NZk02F4y4UWKPz/RUd2+JP5PSCG5avZuD6iSZSjCm3tKqjy40AWHgUKpMrW
pLlI5doz3sGNR1rdqy1bFX4E2xf5JXtSLBayYL0k5lOt8tZYVCSHhmgvcK4tWW6O7RXOzOBuPLbj
yY94Xxa3riIdRbu+pQqu+cOJaM99LGvgxaO6hNykfMcc71Z6QRncZsM5QD4wztvppERtVAQ0EsI4
J3YBNVwfTAjpzZx9VCRUm9frCoroARj3u/6PszCh6BUhYXX1me3RWHoJdGfsh1rHJK1gzOLH93Fs
D1NB16xYsqdV1S8ow0/rWZZ0/4aU50qUuS55ZlaclpqlwA7vCVQDOzl+WNeQvdxZKuAPmaG/6QdK
0EYx+RXmO7XRBSbFqL3awa3bF5XsPyzKxB/xqdUfK9wNjv/5tW4b7YHzEg/kxp0gHN2z/XFR0QWe
jK4wuEnQ3kUQu/hvCxpwVQ63NLGrtQCcGMCU35JGhs1tJF72aIDBkIpc+JUOQU2hOCGcfS734U6n
eagRTeSUa9ap+9tmFQ/NMOuAu4PUeNv5iG8YXlVPIDH2OeIEx9TMh5coXtd4CoJlNqav1hGPc8LB
DAJz0H3/nPN6JLjw9m4K9YbsW+dheeTAd8470OXsGs8+jAs5B0S0a3d9SNKtYlD2nhEEoTCC0Q45
uhco2DJv5FRtUKLMJRxQDJ1yrPhX/8gOr7b1cNcGp8eTOPEXniRWdS0/SJEmAZhwUfBdlOcK5zRW
Ysz6Noyff/dOZtR0xNRRGJ0XK2ulfyDcxpP03S4bMvLIemiNRRLF58DRTxIivG8w4e5ESkwcHe/0
833wg9ixOURBb4XJT3K1af3jOU1hV2ww1/MwMo9VCTi/+BYE6sOrT+jlUerdpySPoFLNsMR1QEDp
e7NGKxHF/BHqqjyi+l1Dyqj+alMUPhEFNVvjFcL66ji73FzG5fHQyWBmhELJ/U9Bkp1aElIVibXZ
CHETg/UTrIRFybUsOZMJz2fTur4Sv89twyJAEBosdCTkJZMsmNexCEjnfPmPBN190m7A37wX6r+3
mwWbX3tw5dYbd0i5FNHFjkEuQ+Qxvv3RmFPVxLMAncC8a15ozFkN/eP5SkG7jsed5pRDUrkO8S1i
g7sOv6japFXqTOl2oOZ81LYDIe4vm56DVYRJPuATJ3BCundXiswRsbnMApzhIZf3179G3AWz/awn
8B3augI5L9iFoeo1BVIoQh4AwBfqUNk+yUbTTkq0lkIXxjijG1kqsdakQzkrdRxCV0lcNVa1OtOd
IaCxvcy4LcprVghS28Gby5bCAnZHCZnui/pTV601ukDtQcGbl8LD5HAeqIDzC5X2a/7z8lPK6tNg
1RmbSBbTpkax4kJVk0h5VkLGIqkZBg6L5AKqiUwHTMnB1kgEKUpaXBevLXXBMCpzwVsjf1Y6e8+2
zz1GptjlTn0pNuCF6XIDuNpi4AXi2eslIccp7Ya6KRZtVDG5GmSyT9J6SLlliD/3eilhZjLUEG8t
7WDt40lorWMzP2Qh1Et19CWX08hpcNAp55EU7zAoK7Xt1OSLq1KW5Yi+Esi7sNWP8wkCM7hWzZwr
awC6eod6XG5/mXyianlUpOoyEJYkjxBOIwRXd0B1B4GQfCuZ2zraqlgjuzpLhvZJgb3Y7gU27k1u
uma3XFqqdgQ0l5GbmkxaUXxmIqOyHU4V6U18AWwjojEPVegmpxWOVEZ7KcZfAoLHnA/WMiSUClIi
9DLl5MpotbIT+Z02BgFLQ46dEhCc+k3KDa5CvkwjowE4DlyAUV5L1Y8UWpqU0yvpwZCqGnD2RTIX
6gyYcxzkHv7hWZKbyauS8wwn7fNm73HH2+QRa8l5ahj2nkbCfOwnHEJMSldoIOR5evd+ketiRBLb
97MOIPv9KZc+2Qe1M3rsbR2xFVi4sizK88K6IUXhMWzPyWyqvC3H9lTO8mivL0yZn4Uq/RjnWSRb
JKQOw+rAVOfiwMP6dU2lg6OgrOeTvHIOpKmF4eZwdtTmbEH+O3NsMRzpJXeT5/RmgMY5D9IrWl1U
pmKdVTrvq9Q/FS9G9LqZPI7ECwlPt8OnJO2QwsBMArtdgNrmeno1WUze4P7Q+j1uKs/0ngl9SDKk
UQ6mbQZVyZlAue8b9Grf5uDFzGbXsHWxnRbQxu7yIUk2X5KxSGoWTjROL6ZduUcvMbgIgmGfZOI+
pgOCg6/WVSYGRmAevXkHQGxOX8lffDqQ7QDUOsmNUNAPzq/HvEhQUKWJWHjWYBMQoXwBjCST/Wm+
SIJiVcImXt10gLSxtULL5RzWM2UOBDESijosz8C8PG0zS2TbrfkcfP/UXm3vP1UAL2DaUhkFZ5tD
PkwQOfMNQj1zPZdVFSppQ4qi/+J4SqZ6m7vW7rFZ0HgLKn03JMQywp/NsZg7ykwd1CX79Fllr7Rd
kLyJ7c3vPFNZ5spL/tIX1OJzfPJGeGTZ/da4P8RRocMI9sEACy+tlclIzwVabsZ2hgnrc56prikc
mxorqBVGo7+5x1b+qKcoMCxVrf1tKLSa4UfggOPSagYf8VLiIIjDmrbNJYa4/WEAemo6EebKOwVW
PPVbQ8XX6Vl1Lcat5tZnxhtCmwTIAsCgRaCpuTVzM7AFsqSFEoZVstoQopdxqR1TD/pacP2H4WsE
QYXjOp2HvTW7KgmkMD2JJNDflgf1JJREudp7GLtxfU/2ZoBxyh2rn+zntbvhIzcFJrzoj0/50I+x
hhjQw6mqdTMn6OYiwqfuQJT5dmw6a8ajHreJG053kX4LS8+ISEdIhYC6vdaINsgDFcLJFm67dti9
LyURQ/yUHdPc/EWVxdjD+c10ZV8ucK+S8eHTCNM75RS7C/KssU7w/7sjTlDcu+eO1oiImoBXt1hk
nZyoQh/AyS1BNN5rLq8iZ+e5zf4RdaSSejO8MdKKQkGqtbEsHBXkpqK89qfCin1GR7kAsN+8Q2nF
NvMR2W83aSHQyUSayumR+yFa8o7tNH2WKrOTe4uc2l/linS2URcyzK4LsbDlUexQYxT1CQ99zg7K
K7OKmZ5qWeYpm54R/k5vi7yj/mA4eHVx7jAz5ChuhUQ3sTgOttDJuw2IZ12pPDC9Wj2cMiQr5yq6
zyFWqou4Me7Gg4bXVGBYpcOoPLTmc4eCQFeRsSQ7NcBHxD3cLpF/9OdH0esPUcTB7mmVfAasiVYB
+5BYSCSP7ygVXi7nkMTu838VPhNV5/lADqyQCWtMCSqZup/x6e0Ewh91T/G79wbWf5m2atq72CLw
l9R4NefTobWkve1Nf/Iztd6evNwS5rDG6WrLB7BIAshjpfZsNUu5Eswzs3/6oBb6NHjqClJPqEqo
EiD4ahLNYusMvmqM5z9+oyOdVvNyJAJGG/6haRKnrAEF2Rlj5AnCimEYgXvaNUx3ey93lv4CD87Q
wBdb2fuO/bSY8joxjGRAYdmCPKImMmHNc6rRx+9vMJtoQ2Gej1Zhp9WvZlWVEVjAk4DN0XZiOGq5
Xg7H5MN1sKytMeSDcjbdgErK3W/HwpoTyqYGE9QPKJcg7gdIvt+cXw3QyYB+xIsRGmx88RexST+Z
1OceOt39RndQOxLF8v0uXxupIjfDL542Z7r/drU/8Slq3yvbX20KcY7Ct2m7FrYTnbuMobrHwi4C
ADfAJrqUBmK+PwrBcUfs4RniWi/GQWSXX3hTAbD9a9g4ZXXRA4ZEpqbQRkwuClx9FO3Wl+rnSZSJ
cSj5baae9GNopXuUITC+C3z+t92diiyLGlLbZgdKowj56WsACOEu3jmWuRTWhNHON7lIbzAbblKm
BidfZyZrd/nek8U8aUVx68oYk9W1I9IKlcNpClUKll/5kyJ86zC7Hv0Z9MyhPXifCMtsIWse4zUl
6w5g75mmceDtxLFJfU8C5dpnCpVdVqhAgr/r5Fqv1QRs2Jq/+O2GJHoVVKuOf64uawiQaZau4SiA
v1uVqd8PPLMIcLM6+8SJWcW61YSu7ucjn9VTVOI+B4g/cV4AlJejptMM4zLdFhkZHv/XzDz9wJwI
X4Oe2MPA7Hc0NZ691eQ8u+5MYANPPI5QMvmQ1A+yLKecGD8ljNH9zWYts37WC9rAgukgTFTVhTpL
4gNGgWq+5mOzDhlV4QrdzmaiPL84BJE1ixwxYhmE5nZjQtcEKelJClFOupyZ5FqdyA06P8GM4rPH
AOw75WZvG/DtClfrpLE2IQiWIiAcQ03T7SsUwbf3gHivxvXM1xJrqXRRUeOR7ROPvW2caL4GERru
UFnZ1f9eq3Uhgcsg5McU3bY6Ulh+Avr4kt3yGvTF19moB2gB4PAzVF81lG4T0JSpQjPUAk+nU/pO
OBvHrOea0gBxmoqswSk9dEvWN+RiKABCL3gL7dMyUZSzOaS0679I9ll9J8Vu71ZHxO5SEAna3LSn
WePUX//XIgkD/0Zp+lM3iIUnqiqhOMr3fnH1lJ2tZxGcxYnjj30fJo9AnnawgcKxvd5QCYz8S7W4
f430Rdb8zq8ezq0YyA8hI55PUE+VOVKtlzFLuHazisaVLw6XkmBlheiL3Vz6SGUUUAQ6IyZiNwiW
VDLE8K408PC2hylUWm/X3G+fue6c4mdYJuhdIphzSf9MXfZ3GFbAd0V9pQUJ6+yj2n8WHb/CEI3T
nH6QhGHsa+uJlTj4beH1uM4/c5sK2iSgB/ObFzVckQaKwiP7edHgtvKRS5oBkpaQ6ZkHZSK4xoM5
bQT683f/cDaZS9590a75lK1B6tbpfVoQ2Io0x17ca8ELSwZb0tQ7NDFb0KqRYvDIIc3PYjQHLmu0
5u+li8DVhWIGmpexMpPmsASZOUZR9p/B5PLXSirwIcFdq2Kh2cejBBXQhjmOgnneY7FOgvm0LY0t
+Ntyow5CFyzNWLTrnNIuTv8u6tEMAnnCMPEglZPh5d3/jjnnoUX85pgiCPdTC33lYmeBqz7diEg+
Uzuh7NyPe5OQ1yT82dDisZlxym7TDe55G46yaTkOkycAG24i952WFeJiMlQMu447iz/RgZtt0fDH
fIKe7WJovANwzEZKut5fmDWFuizFUc5ALc17E/54ib2uteIbgIjmqJSKz8vh3RzpzfcDd7xn/MR6
vGTknBC2basYexIA+H2oymTARIYY15yFKZe1oKjaVengTW5zQa1V7ooZR9FePDbPbzkJeVlKKrZF
fpY/nOXmmto5MFvZCz0f3O391hpwEw3zvNE4ipbPYyGseSGoUGcRR785SxxAP3nZ7fHKMqfY20ZH
6usdYoRfvc962g1/5N0AHPVM6UT2CbG0xI9JnR8erhtsLSX9jjkm7iC6leZDJ3wSeP0icwI62cH3
FffocNLB74cQZYtg8MK0poXXVGC4Gwtp8JZHHMGPlcYMrpO8TXtEkAaKpvCzTN7WvlHC+aLoU++T
0VtyUAlBGgcl3Yhipf6KuoRfvSROdzqySwEvf8JSS+22iEVqiVZCGtnGQO3nWiixI7XjY5OsgeWo
8VzhTavztkTFikTrtRap+vfOUdzlVGYCyorb7KxbUsDcyIPiX44qGDS5HzOiClBYyBl55+qhlATI
Wxd3NPrFwrcNP8d+XdkP7LSnYkMPoo0M1A1YZd4gsgzCCnyZyXBOLM5/bGiz9ErGfGM5mt7/1/ai
ck5dATAv1mjEuSlektnx2EBQ6weYpKZSkWchMXLPrYs37KOh1HUGLTH6hsFKkjnZeUJJBb8VFofH
JzBB/MrouAWa/bWJ0YiIuXzDgs8ce9yaxI+tztqbhWswjxlD2FANUEo/tvCXCZ0eZQ4iuCoNmFju
9cIW1TmIuv6ng9bcConYEv3A1Ui15SnYw755s03P35/uwVzabXxBSJtjAOJ6M+yMV41Dcqn1ehxj
zEdbWvbbafnxBOuxlQC7ckQAKj4GCGl9NpzZq2bILE2u+e6GWiPl+B69A100jQs2tmyH6kfiCNbO
o7/00PmQn+kjYDqWbvdBSY44Rc7LfFjqNT+FrmH99nvJvo1/i4r44X5q+v5w5XbqMWuqeAR0ysoa
08ZZ1y09Iy3w79Qkxq4dPwfqA4jiDbB/Jm43yq+dNv5r0D4gi8aCr/aRnZ7jgzqxua89BlBQJcpS
HlxejTLfuqYgCCBvyKTYVl/hbXCU6DI+pc8qGjKTKRAmyZMaU+5lKb06G3FkDbiGCbxEDrxjMjZx
Nq5IyaIKw55WMbEPK3Jm/c9QQIPD4r6uBQLNUVqN06IofFSLrT/FkRY+FA9ERc48j9N5GVIa6UNL
oxSR8e2Me5XVx1ipgY/7tDPoTn6dkw8nlNtgBqFYGMTloWmszzlQ9Df0Uoz1ps3jq9S4daRTVPUY
b+qTOLAW5oFUtGTz97yi9fKTLd/ZlSKqSuNAgTNe9QXhjmXi+v8fDW1bH/KTu6+++c6Uq/P98JJb
hf7QvlMEcbmLmopiDHjGLL4plXmcz0quV1E6/LNo61FN3gaNBUBFhjOUYi4A6rbGOR3snTrE+4zQ
o5tpSvH45ELDtaoY30+aALQYBd5dO3MneY9gRJWpRcPfWshUS0wHqlU5tQGpEceqtmZz7dkH9TTw
HmYJW6N1/PRFHGjxWz0X5kBGQbngl5MYqinrCTtkYdWALLnFpb6/2WfhdbMr/gHhU1gkKdsbNVlp
uC1a9+oeSAHYvm6FyFFvNK+flxu7pssempWBJc1NlDHFF9sHyb+xEtyR4ZPHMi5JtkreZrRAkIip
6vADgzynuiWf8462lJjZ/VgAU0LUpV8jFjKYu3tYVnr/OVK0e7FQi+PcsV1R4EOq0czQpKeB4nhQ
j5OT9gxX9w36ewOaQgxbLqxMp0gZqtkWI9ngY+gH1vzLGq1gAmo+Pgms/37wVdT39JydMlHBmNKj
NUURxmAhrH3aJyMFgpshFyN22QD4Y+RbKzNdPx1uLKqUmcXLESZMQ6rSBVJA4547kFC0MXQL89gz
XuCRoU9l87YlFvefFYnR2G+sB49DYKhXPk8IvHWXB7EmoezySSBuOWKll4IUMOwpsEwexBISJG0h
0QeSPaOPhw6rDCls0JR9myZHp+i2wr1QZbx6TVo+e+9T9pxSOYznmdjK1PxSG18GbyQ7sxHLdCvB
FjlL1WZbOxPc7L1tiFZmJK1rh6jvWVS9JSnqUY5iM4P+nwaMjFtEWXYqCBf1sppu+R6nbic3GaTI
u33paECHka6G4Aws4ARlzz9hRvcCye/8k3wXy7SUYCE8lZBBAH1EE4IqkA8C/Up7h67nqTrVKIKS
PYKz8Jvs7bp12GQwiVubeYI20IDXqZRNuvah1EzlZw11oMxlhMuPAwArJVj3bs3+bbj2RqqAUV0V
cLvUOvREmV9ucjjhWDNKeD8jqAz8OOQ5qHVjUhx6bZGAz+1SyElfalj5Lx9JcrmOpzYKXQ5rBAQy
7UQnEEcl1sYRhpq/97PwPvB9yDhM5nfMCjwBnEW/MrHNyyqDqhx9g//AvZSLkli4qeB7ave2Ff0k
czQpmw0sZeYlXWfAqqVY0SPIPJb0DUC2pqNtnineuYvu8FGjmEWDmKPR+yylZcCz/9I3YQOlkSGD
oxv7DiEWpX+sHBCg/oW12lDa5Dw7lsJZH4VeI9arXMnr7yLAfPCP2n6MRPBD08GcL7Ss0Ckdfle9
qgD9NDNy0ZqX/08HgNpildtiwlVdVXWvMTg52XIPJtH2eyUPn6vF1mrgxjKUrO+vHa7RD6oTp43V
kUKmc1FMUChvCIbooNgkFEP+jCnXnO9P+To9XzjoLntg7n1GuLkWyI/cvMMSdjukx7ygrsL9lBRA
9T31c3MBDqaUBhEi5Vk6sCcsDc98iRfaqeBxodtFFlhz8hMni2dtTS7hkwMv2mqulpmP7jmWq4qy
srlz3i0GKfMqz1MukFhvWitt3+rFRm8iiGA8vbsz7zMgeXZrwDm7YjEz5FaIQ81/d9WGjd7r0l/S
0S1Dz4w1hycqLTItiL5wgVsEPlXsPz1/FHScF+z3OmI3dV5WifEo3oK5cx3uKH/xWLQ1dq/w8UTJ
wOBt6ZOQviftv3PzLWNe5qoVkrL+idffDcoSFz3OIOb9CVZO/p9NS1OpSvqcb2EjVqi/tlnccBNh
TBgEJ8p9aB0pTRxEnb0StyII41vFhZrcnhz92Vf26wt7T+/3RIYAfcwLJs5ng/LV20xHOoEvNIQG
SFNnSuCqlfpOK3PZQ4gWgoJMIzthb6wuclAD3FUFJ4BQ9EEfkWp/93UuvmqpAEBcuLBnPTXISfFo
sX3ueizqy7y/GsL+IwOBapEmHVa/Op2wVNRFnI+w7AqUFoIdcTtIz0mY24EIc0wOfZZ57zelh2aF
ut9HvW3MiUQSnlFLp/pdQ9nUk1wgJU0conFxLGZHFkAbwzKGcGdsEUAT75Gh58huW4mIzHX00Zul
0zfY8dU4IoSiyPzi5mo1OuN4xJHJ3SjRuKh0SdTVJhsHZ1YREaT3Lc1xzTrVxC6ZeR2oUcodAxCd
jDe03z/8kMlSX1wVqGGNq0yLWcI32t5GI4Yrqy1peDhfFmie1q6EVrqV41d31aWBZRz353jJGB6l
hW0jTJcSQe/GED/qHyNf/AEHVSbzhFN0j3u1IvEvzdRO7YQutW23aytGJG7iOrBkfg6brs+ajFhv
GirGBxvyL5yYCniJd3ESYFfT3MXwGVqcUaCNufL9D3Db4/nIEE4MGaLMKxtjh7PttCJTsKoI6tm0
TisC3Ss1ZcFNkmY8j2OMtSUH3LsPgjeij/D/usI3FXpyqEJht2sTMAD4UvKSPvu+bV1eEcO5IZPo
mpgO3xW9HKRIyrvQakJn1XY3pFXZuXkZDsBr4/sNzTS9qIRbDdz2VgEHlNC/wnAYt9gTXwMQQOKF
uPoLTYjzIz6KGmgCDHPAJ6vkYbH7DMX4rtiz70XClsf1taFztzkKcUgllD17XH6oK/9twZ8cbhJm
Axl29sRDiYY9B/yu04lhn1aa23nfHWkxrGPRocgGmj2Xd/7vioP971OGKIKW8dCXNYuOlOFQt20C
p7uOH9vKRT9HtfyePRW1FNQ3ZMjvPxHOUFyGlSTPt7y44+57VBgCpxAGCy16XcSKomsy7kxu7hFq
LWWgP/JIUAn77lyo8qJTDpQRzIRbQLWtDwz1jPqZXWCIWQhaEehhw9IMszQDAlxG2XzWBz/Y4zRI
UF6xGlCltcb7/L2dO9NISAoZq7Uw7hwc7qvBxUQFPr9OjUfd7vIPu/4fr5XdFT1ju7dN2xAy6zaN
bnZRiAAVlAnWJdkqT5WaId2r1ebVZjuSM/NMoWBGoGd25JzEwCBfXsiJqZiWUcUUpsooPLlYgVCH
I69+3TxsTphlal7OPwiFfLbdfvXpsi/1sqY/1x3dWdPbwrVG0dOW4AHhJNvYSscqMtejBhLV1oly
B4hpVQ+i/ykYLOuJHsy3L35ErhNGs0BNdEOknepXWk/m6hJPxzUh6nHMKp0rwF+JGGQTt9jd1prt
AoxKksnAOW97fBFCJBt6DeSEMjPSSJbum0Q0BXb0HQLkfONxO4k8b24PKTEblYiX2cfJo6VTGmQQ
DmVJAbNyeL+JsNjIUXHepsT5myrIyfEpHW8ukSMRI7yvVN6AYH1FmHGapzMAAmRTCpTt84iTTRSk
dT4YbT+ezfQ+CZk1wj/mZ/F3Vu24N0EnBScpnIVgovRjedrXFsCzFzs2W6XxCoXBLMAtOa+qwysd
KAI5o+9K/hts5r/mRwywOiX+lLJPln0EIwr9lLABURwMCeGR2hXtajc2wOC9BojN8lQTZRqEF8pe
YYMXd9dusx49oNCyyoxABjHbElNanEFUFdwJHDphVdviKxnnDJusiOV1/1F0kEBb/WK3kbBWn//p
64PqAxz/0DoG8tCLAilHqoGxzS5CxjchOAb0oQSBGOjvn8dClcZQjowQKsONPJljNecF+jCJYYkE
j/yMqF9GaBfVuzfBHEccYlbTH6Rn2u5G0g2vnJFvaBUMqIRoJTQL6RyxHP+RMc9XdpVKTbQaDhOH
UCRwyolI35ycH38NLxn4VhHUQCavkHRsovGxHaqBljPfGTymzp6NlX3g94T+aYxxr22Whq70RplS
fsQizEO1AcbtrHHOtxsV6uGrfQpy4eAVnexVZSncZT+KzSW8peDrAsmrEXXZxDkU/FvZW9DyuDAi
GWLIMFBiXSAlvX5UpkWxSon8GmkFat1RTH4+W8ivkrBXiEi0m1Je9jo4Y/7m6+BPSdhL0p6ZOWTP
d2DtNlT2ARc1y8sHZV3v5L6Nllw8mwBR21daSAT7QSZTfecPW+x0M4Qn+w+VNwQNSJ2CPq4RijLX
g112XVa+neygKhv60AS4MK1YfmdG4psGjsS7yDfqCPIyhSL/ronGxeMzlv1WzT82fcAaxrf85Wov
HK+MlGGOiL3Ci7o5deJ5P+xmteo4KJBC4CPb+cYX07/0Zvhn1LKX3X3c9ghfXcRFTgnDpYIsIYx2
+L2BJVLmLIg+g1uKOyvIItUOZfblWHp/kmytN8luP0JjLymfTbCi0ttLUwitkYD5YEeVtXJ27aWu
Jrk1bZ5CUiWidOidEwN7OcKMrdUP4h+2Vu2omHrbD6C88Xoppwk9VmAIEhk54zJVMUuIulyVCyYB
GyTFsiN2p/f1lRvRsWs5cvffPMKKm8hLwiTOK01pFs0H07cUJpldTshq51W3xyRGzHUo6K4xqv/M
GKb1max1Bb3cSqc2OhrOfZe8nC9vrkKjFRUFm2nnHDxfLgJ/ZtZTbwkG2EHbxcsbAU/UzAc8aVv9
JmkiwCGUSuKlpy01AujDLJeS2y9N36hp4pAcVmL8msiMDssynEnbep5ftYFHrf55PsNUWHIeJfYs
hlytpSHjnNfsGLAi/pH0pWmunNnqmT3P9/+9CQcloElXXcA3Wz+3UjWj/Ss/tIRhWXgo5qyB2CYn
HZq2VQX5P5JefrDKwoCTft2h43Llvq9+uZZBNx0oK+9Y4uCeLuMyjByIuaU3NgFipTIA94DLSaZE
N9+991i32hzSBdp6r1exVIBgKFUk1z2S5z6bUdetFRAEsIIZR/2b/xAf2VtWm2v3XaGWuksOUnRG
dLuqv0we1yfuJ50a0dgbyns8oAv/XTRLbmSuawGo73c2bl3T+28ChcSkl2yVdJAh3OiSWMkSKsBy
9vgAqhZHsOq3+v2Piz3N2BaRjdu6J6YLRxyPzmQMnoLkTtoayHeTVv5TboHW7/1sDt5D4ZTIcylv
mhs8iVq4Z+j3TVS1uSoW0kIKMBxRrUc4GBR7TsuUywGmbC5HaRZDqgcpiiqF37GnsEBSUIeRcxlL
s6/CS93p0d1ybuR6clA43ASX/Sv9Lbyi0KrH9X/IY49W7eX69tvVCTXlS26NQOt4/QahpIOtsvF8
ft4hAD2EypQ40S+GVh0iOEl/DK+T93IWP1JiD8iVTn/JUZft33iKLGu8YM+Qop0KF/a6dR6x7hVX
w+ZZdUa3uGeUjncroc256MYI53w865IpnjmeLRT1dVQiPc+8tFdf7ZTM9X52oVLkczL9q11myKlh
rBjQwxo2ChaWZPhBz4WN8AY1AiWCKEA7jgB/fJyrybgH0VMNZ88fTQKGtU5liS+6cJifMLilfGUn
odbku0n8lh2jC1Yvu/+SaNUmtOzxGzflltOv3AjtdxqWKSidPvjFtS8G+6kG+dRNFZv+60wMNhKg
xHn5Q301QC1qO7rWpNWjDClqNacsUbuoSS6edVddAVUc/MEiUCZfockf+Gc90dEKH+M4ofWFKXNH
IFKS8WWBlpznKgnk7lIxNGwOMogpw8xMdfZBMf6Jnw5P0whU+zjg/crvHL+rCcyuR18wvl02a+ZF
tqEmKnXr1Oz1U7/UIn56pMgcPJrNHShvZPVnmOv9gefrxRnPTRLehpXWbwzIERkwDOO5hjne0YRL
MyW4j9IxD6B9tv88To6Qayw5/LHN0T4M90kecoYhbENgI4R3HcWXblzlH1TR77fSHEmL8j9233/Z
wT4SnhFG+KJzNpIR7HS65+eUUyVVNMwo2EfLXjNEvTVXdfVTEnlLLyKORf9hJF17OMtRr69MecWm
LIjBxCYAggEKK8pdrspsTStOWt3fR3iUjgU9bQ6cPcOJm1f2ZTHjw1bnPhxxxb8TBUnEeDLqWP+J
qwdDAShhr3sLuUaGHPiLY639XI4R7i/eyZPyHbQbHed/uyycZni1qRimXOMvMTC9fx5czkp9fS8a
4FjrJ4il2S58haYxzbkfjDojnPNPe2W2UskZrKZ53v/00WenJLC7tRXsQmbxiKKU31baQ203ue6H
wCBECwhtXqDR5SuibJuCAryrtHz/GWBZoxuVimzY6sNZoh2yy20isVL4/rOFkQV6obWAXswZZEUI
3QysOv49CUCPZrmycnTZb09mLRX2yqYVm4abGzx8pgraqJr5w5hOB/fyyS9wJhvg9f8E46/JZfoO
BwjjP24nrzEge9+neDWlefVTjq3neB6QH8f43xmiwW311UPYBThQ1barvuxq9ymIE0ZNWQrM9+ob
ME4rH+2JNMQVyAWidELFIBi0eJ/YWTx/cTY0YjYRK9bVnH6mvf4kbKX+B9IKSnYFJiuI9y4UaPpx
PxryqP/5sqFoYh+jitCHVaiF66g/ZBQr/3bO3MXrA8Vy35PgN3aZBJ9C4yeEjoRDx6RVBkmD0VXq
6lQKfx47CtchTjgOU6EnECaRG021rkmMmwV58237svoEJmHOB8HnQ1iiCcwtRvCjMJuywp5sdwKG
sXzrgF4s2+bQFT7ztFE1nEMoTUWY8ZSi98P9Wv9u7qQ5yY4LdOKqd46uzZYciDbwPbMZMpVyOlZp
uDaECahsib7BD/McJ9G5qnSCZ5MPmphjx+JoMuN+0efvUlrdHxoozjA5/Cj9TlRkccaFNb//vJBS
g6P/JmMsTl++SWu+zIbbgCh5xLV3hM9w3TGNa18ZVYLOv8n7RvayQFiS5ZC8CizJtc3CzxoRSyXA
+JTDs2JVX2HnEczDvU8hbXSJHEsBux/Qf+3iHJhq8RSuyCVGIh8J7WhrxTdAaRpQenXB4nMZPNh1
HX1PRbiKDh0cd2P7gn8eq9a5UembzSaPMJkVbzHgTpPw3apoS2Bbwo1zocAgSMuU4K8OhGC6oftT
7u46T+UrwIZuvZcgslYniTJIxTLTS0bwLQv9dB4u9D6D+ubagL4eSRYVwasnnkKpNY1b5XD+axmp
IBXNZgl04mctQo4OIINfL3T2/B9W+E79fO86cRDtkhTTFoxVZvkbouelRhcY1/koqXLkOYmFsl/f
rlSrvwkLJ4ibv6YtV2Nq8yldfFmUzcgV3x3FBARvwFpIrPUa+Byb/3dbdWF1wg0etC1i6lT6NPf+
qH9x3khC6xNceCqP1yxLFo0qIup/0a2t5eQbvaRReFB18F50YLHBRHgkh/i00YxtQEs3vH9FBonk
xS4zwRK9IGDtUEhJaobyyEyFiBkkcuUm8u8+pu0sbajWdtLjCePwvMqPasd7XiEYLlrM6lwigv8j
wZa3bYkeMc4dF7egtjw3ej4ks/56kUrPgbzz+qU623C4UoIdkBxd+3IE4Elq1NcZh33dBzyFqEKL
BoJveQYwhW0rtIxuZmFtTCxkrFVJJrSoaDAIrlqNuQxQZBdDkIzbAsi+38jMa0qCgN5HpHKUZm3r
IPwkFnN/8guJxLGkoULaKHoci220jlqo2uB8q8aRvo2UwQ6qWyYyLA/lXGmetAte3BT/+105Rk48
+v4T/aDlAJE3YdjkjTa5rBW+fCGLEYCUUHHOZYqfI2Zunm06QDJ/mmjB6WYoYkHTYyWs64fSOUIB
JWCG89JrG/iz+48L+D/sJHWbnsstCqstngscKYia3/cCyIEwxkTsCt9EEMy8pmC95WHQvsVX3qfe
UxRQ2eWWbWCKY6TsOIMZq/kOeRMxHI51/dPl/pp8A+FqhcCAL/yDTMivY0fpWkSYNC220xFG3Flc
ZZwd2C/MkpvBg7Ip/+B5NsbzGqe6huN8Yv2CooP/fhfUcH1axvYk8nQl9Th/OvZVQAer9ca094WH
lXqJblw/uiNnUPVMHO5IavfsCV849xc0MrZby17dPdoVntpj8LSgVO/Rj4wpza2MZAWeCtv5Uoh4
HaqpEZLkPnDmpkptO4rr9451Kqbs2T7HB4lRNRP76MlEYVqa0o2erPU9O3P0w89ul0SlY/tYFDFl
f6xDHuvJkI1BZIFU0Q3IU7IK3ebhiyDpNQv42HzDzv+aJjeaDVYupytsdYXrpgJaMeJZchrli4ZX
6JywhwKFps81LcWnIpCviJz5q3vqUk6l2uw2oNKYL7gNKkdwoQUr2MIxupn/gPTfQ1DJ0EaejyRA
WyQ6aD0ZKag3gc498tpqcq8ilBhqt4pbg+ve15ZNZco8XfCwE6nKYz/e84kqp3JQIdRXEh0PLQDP
3R9O5QE2vmvOu0ZPEUJZ/DPApPPxhbGf0DfAuukjiQw3hX6o6A2GgYtBFDaurLDYvf5oE7xV2eep
gmjB91r8MGaePb+M4vOw3DRuGqhmCwFluQE8K0rB2m8yZkv/FC7WhRv/qNz0pf4opLNJjFA1ASST
gA04OIXD+vuNew3Ucdafw5DGfLoEvbgNKN8FyO4xTMo63fVQJwwxvNhwKKdWw08NgiCY5nWUiwwE
DsNjk4RKcLgCdi4C19+mmnV7G20lWo7ikTNYtoK7pyvGWAGzpMJ8XicQIGRTjlBNRxnRPG/h6RBt
u84m7QkFy/x3mPo5C0JM76Eub2D/IQl7NIOYRGoffWovegTnGEZHJThVJGDe1+JzFgkUJrwhEzX2
poU9i+wmqivAbSKMWu4XnObHJi5wZwNhK4neZskPBGPyDqKxu3eDs0as2dATVFN2uNNdwHtjtyY7
tfMqAfW828HFyPLdfO/4u9ygmnXcJhgwJxp8SBy2lG1Uw64+5eZsPUECHRfwn0UgONjSjPvMGYd9
vlKTiCONseBRskBdz6+5Ixi9ZhMsu6doKB49slURZ2n2Tl+J1gr2tSdGFAbI0HtoCgT3C7sDMaxb
mftfa2ndMop1rbKnZucolUx7UY8GpKcbQPPGv33s/VLtIgxKbQ5PvbxhP4PJeh62CfAtsJJUlCkz
TEBjS9B7xpV12hz9OWE6fBayVT2YeRX2us4QywrXXvX3VklGIu3R4AhPOP8JgMSe/cIh52F4qZ72
qD9wfgLz0xg/Lge90AC7ejlBd5sS0fi4ftPGC8eCvTP0lgNZyJrGSu8MEBogBnVOUbMDkR8+4f4f
AdvGhiTyLftQdzVbWBB0HsxZ2ZW0HTo3hAnURlfJ6kENM80e2sQoPfmq02eItHpJBYQ6z1yy8XmZ
Da4yUP+ST/Ru2qI53FJQl+pmD6xzM11M8Ef0u/jClGWw3dOW1/vE3Jx8gYWf9UIGjXgSShuDpu67
uys1wgow1DJHfb7bGyEMwK7b5dZ81fUcmuqd1u4l6PowC/Guq7lE3VvcOjfHq7rSw/DIC/+OgJv3
3R60FyVeWFC/tB/mH1MS3wFxb+jKzv5E/M5FRwmcUNfZAAamU1vCT26wJs/A0ksPMQzN1FFpTpKP
kbiBpjSojjmtuD1uoM0ca1YfH15Ax2XPqMPS1xRPCYfUN+wziYD6WntGlO+CxKIAFLxAuX9HvMBX
oMya8IwbrT2rglEnn3EcyPJc1ww/r//4cw79uiLeepVT1WIXBhKcicsb5pYVVRJi4YlCILdQWFRX
EFYf2cywtrJ25a3NJp9TynKzZkODhdlQY+ShcB47rOwhhxfCCEmxnv11QWD9A1WzYM+wUyZnJ6i9
Nbd/W5EkihhjH72pfwxt9FtY0A3XCyZWS+wzj/K05CTDZjOyDU03LdQQhGsaHlvVyrnqZPOCYoCm
PmCo7Scfobf2Y9n5oaYrs2s/S060u4mtzYVjhTe1gmTkoh9VKGbHVtz/UGz9DoT3TY1skrUm8mBw
idqB3vlLkreV+9YvaPjwSHMlRDVSzPbmZ5mwUz1SOL6kvBwp+Zpg9GvresgrSTgb98ciKvxLGkYO
tvw0AnNHE6rUy2HBY3wtxBFLUw5qkSY6rsn7DlJGK6bb04oaYoUReVIuJhT4o/7JMVvXSrC1U5xA
AtSTVxNf73ai0jXel5OobcaxUpPHKwBTtCNMVeHwtVlRM8FTJZJKJoDCc/O+IDDPLYTvoE2DuhJF
rCugqKqp3W3c7oQDhjOWGBQaj00bckzpuhx0odxg5ijNdiJHCt/S5AFN1PP0nsPE5H300FadsnFn
lHkGXQBwdUWfH2uandFPyLlss78TX6oRFo1R5xEqqSJ81bDr899c6JWWIRFdgStIfLRKCEyZySLj
JmMg8IyZdUEIKAuBH8P0hjHwbJ1bHIYOiVbQfa46WUVTL9x6pO3b9s2S/lhAiUU0QuWbhSj2TLvs
+S8+TMgWo4PacAp2+90UIdkjO7dHtHKoW7xtzokeJRNo8Ft38X15iPNKxTrBKtSJMeZWiknWWiLm
3RWzuD7pOHZGlW9quCeM7/2XfnOrlgo85YtVdhJLG/6/C/+8vyZ0/vmqT89FKfGzw0etzCm74tUW
mlVZgIr+oC2J7Kwzefaa0zMVtJsq/SbKaMMRtjw/GTcKoPv+Of8KVsqezd6rQmSHx4ryzQDzrwIk
LNJA3fBJ5e3eaSMjbmLmt7lAaQ5C6XaktEcl/SDqMngHTIkhFaYpw3TZ1xx5EaXUViBoR1nE0BvC
5feMXL8/88W9tjGlrYe72UiEOT8WdvTNI46ani26VspqUFaUEUI6rrixMIprV++3Oiw06KjOKKH/
4AOY3g6GiRNv0Y3NaxR1rQSHhmKxuE0IDd4vhNp7d1fsyJVyaqO140S/1j8wNpCb8nDgh1lhDYWY
vgFqGo8mu/iiNaCssDghj7MUxwurRo2wljioK653pKK536xhewHjgNDnfZa3r03EAI04Nz3yGmsa
8ot9UVACHCa3VXyTNMXQ6kAlLBoWRWpwK9294VQug07fzHg/1qSZ7rEBBPuPWeoFP4lYNhBT0Z+l
Muqo95+hzSi3veFM9Q4ckobEuJqcHql4DFqo4VsB8Q3q5b0NZje3B4LdUSmbtag3813Sr3H9iCyI
ok18d8E9mWRCQfYWcWr6nh4fYUoAQwSVbzdGutW43lb4Zb/+qpaCjPUx2w93WDwfozSrq4BdBIoA
TOqmd5n6tFFmxAofr5T8HJDqimynFoKzl9RyolOPQmi+bBrBgO8kTk7bIKhQ2VDAgnmFeHV7cj1f
UNtyXeMpznc+rAL1Ru98i31HY02YuUSdVVV6NdMiIZTEQGc45xCiul7c3Eu+IoDWnMW+Ukiw+KG8
Q/Ow75E+m1f7+XN2iTSQJsrNeax0QdiU1yH0RUMNJop2hoWYT4HxkPa5iWcNOr+rIK4cwFMBPDlT
+LFYXzeMu8DMANAm2tZSyfjVLItEPQ7vOIIe5vpdGbBmrLh3kCKcQAYh7Jg9TuMDUXfL0HmVRBlC
2T/jQ4mL3rHDcRAITnJ6/gM0sosYzYEYUCsf/voukCsBq3jpPrieuvY8bzsV9QOaPs2/8/DflN0+
hqwu6T56Uj/j8WYGW99V2ajX2n+hU/XZbhIDYs/xd99L1HBMGIM6GnkDoa9nOUA/ux/TsEKstAMJ
uDHn+13E5kH6MCvakE25QjcLankEY7s1nfBU/yh8tk0Hhtth5+8aZurrjyYVGTPWXlQ6Ygqo92vA
ip2ZzZgqPZdBVYNGp9lUtgESHzbLK4q7za2vlmkZbfxbgi+0BPYoj80KRHdjYY28IBgkU79cjTBq
S3zG0LKTgyLiIexixg7w5QPNfCZsXbV9wkiF3CrN4KzvH5T5pURqXocwh4xr5yKbwY0sEtsqxfSU
NwjSsydVyuc1BoRYqAdetjGC4eB3MLc73j1hshjSnsK5IeEE4uFMp+tozmhRaGD46HF9644MiAVY
dMti0cQF17e1VKCoWSFRK3Tky62R6Uok6jbk7ebldZi4I006oOVyIUqF/zhPjkL0BhJW7LXFXMk3
25qKQ9rXoMYW40WdSHVlqt/Sp0QR1kCz+hwiUhL8Gv9JGBolaz96t5Ni2D2MDphh5QZTaHmhiQlF
Tjcsfhr2I75g6tfEXPoTuHNeV0mFCWM63X9WWamUhtz3WtK2mJ/BrkjzDGlJG110v39PI8fqj5W5
0ueOw9QfBk5VwbZlRUjzKazNPnf/DjKM9etnb1V3LSMydenLBuTPkFlQeiNXBPNRAOsTWbiSoEXD
VkmvhBbzdCzJ+kcVE+C2M8answDYaTQSvjF/rPMdP2hxGdyoywAMCjxQbV4vY9oH/0CpOlfUvbp1
AIodhkpb6ibH+Ylyez+T5TSHypE/9W7AoNoE0I2SH4uoXfS990TRxoM6xt4+0MfHEUdE3alf0XN5
eCamqHD/Y/JVm45kxY6/0xwx7HImCBHkB8ERaIZg5If8vnKdXvuVt9rnQ56pvFuLWyfkr9YDPpEe
gnUnD4iVWX6xM1LavlFR3jID72JXmOSIS3zl05vbpx4Kg8bAKKm1s8dbttMBQw7Ts88KXuydWObJ
miScGZ0do6T1R3hg9sOm1KAOcM1x1GHpMsK5KKnP+As8P2o8IoveRADsksnP0uS/PYz/ZTjbn7MW
OAozOmN4GRqAKuXri9fOK+IC++yf9OFJ01Do958799dDSEJq5KAeqHEtvK65gXhU3WlQ/wkCqoWa
wSoCSj5TZ3mIz45/VC3yYtMJzHUl1tnn1QOjSq0sWH5acBfDnv4luBhNx6t8524QqJJRt5RBUR22
IA7/gifMSlsKg4CDWSFLHjHDvHecXJgkftdcEJdb8H7Wg7Gf8PhnixF9XHWZOCnMGfQDnP/V0L9j
HnUEMt9rA249v9v5HlZBP2qlu4SbZBUTw8H0Wu+u3QRwvU48DlH7tn58u2UgJMrnDlMydkSmgej+
a/1gpgiioedAOWmFF9HaaW8mLNxJnYQ1e/1zkrCR1pKcTi3clO+pDcYCXnOblzgc+ver/FAG/Sil
HIMXywX5FTVzmuS/oq/gbvvVPqd3KUFAimCnuXlGm0fMoqb6Z2RaRHg3X5KA1neP/bzRqtJ6hnXc
w6jKah1WVvsHaOkQzd950XVkLX0MfWxZBp4XRENC1AtRFgPtIKLtdV6sV4LpIcATFslakb0DEGcL
c39XYqwk1GeR++xq70E8WZtWT1mTVO/56ggmI9tgfEdruHglVfJKud2TBIFbo8leXg/Vcw0AmZof
ahRq1PmgFbvPVUeHJVAOnRr0Acwscl1vYxF5pMT+k05OVMLEqZhMAG2ZYZ9q2Ska79x5MWI2UGsi
hfvuWU21uY9uh0D9KhWFWnT6D7Tl8w2qYdRDFcr7e/RUIw8MAInoDgjiAt31uHN2jmjo9yFyCjRS
IM4apGkf6uGqjiZ2bb6ZnNmwtC9II8FBf8a/NnukkPAAqQZgMURa4vqSPW8QsTbLLWB6cCz7NPDe
fw+7K+AavXR6ROquy0+/qDT0ZZo+7w9wwJFEhPMvQq0wsGUGXLv7zk0+uy5ZzcuE9gscQdIEc8mQ
vrWSGNeXlaAJWLKhjtsmHVbnMLvsXxviXrjA/KD5X2lgS+UnAvlhg/6FKgxjjlDs0wDsQ8ZSqzEP
jdktxUQ54OrfRTjJD3t4KYjAj4fhpJwJ1q6fPW6v1hgqCjdhC2V8Q9+l82FOFf/xDAAGfY3KUk6B
AcOP/ixhjBKnVUEFjO0StcteV0moWHltKZ2rvQyrk7gfYDIli9X3OixKJQmmTVR4c16lWiCSspcA
y3X/MYKnPWEBZrgAqsGl9J5NM5u+Nskh7kT6JiRpMjUjGqBVuHVKt/NnJJE3DHlUo7yGXrAnwxR9
ch4kLUpai172+a18KjK9gkndtXotSD9H1afdYotllOi4DZsQI6FfMESq9OeLoGiNizNP95Z3plM6
fhDvmp5BvrK+e2Nqca1Inm8FZvUXD1aBOUqXnXDG6eflgKK/gfaZslj/DRIXdga+X2289YpdLQPe
Zqr0ZYQla56UkifP//Xf+FUPjtzomNTVqQpqaJ597w4grNiGuzaoX8rPHca5KaFVWO9QLFDEK0OE
SiVblipSJsQJcGRJE7kBWJaP1CEM9oJZRJMFmhHd6Tx+7bhPBQ2sDwCOGxuk9kx4RmYFn3dHN5C7
ZOTm+M1kjrvMP2LHHMeOxHRnbhXfLUEHJ0Ny6ZcVFfw9noldJYOtOvfAdV8iGeZAXjfhS0ZQNxBa
J+BWBvvRWI2Gsl/UgBI2xrv8VfaC9eECs9prm8NH6Evp9XQdbLZJ39BuJsvJL1K5QImfCFjhtLOA
P1IVn2+QuyUy5CJ2P1H9OnIXd8DpvPX6+oeby3+6PtdtREsZRzmekxzKz7vrqCUwTN8iua4o1FNW
+dOwmx0gGwuPQpYGwp2e9qlhRcawkesq7w1cvEfjST0CqLHqka7L4xdbNbYlIsBCYDa6JahpC+7n
LLe4o8Eg1r2eyHEOQeZ2dSGjO86WCOG932u/gbvD4NvdBGcgQqlyNh1kfKK6Taoljli8/CAkvfbj
jb39p/nvWjzGwZlt5AmIrEG0z+ZcwxN9VSuRnSDjDkstQqvVANMzueh8+RM73UPHCpbuMV6HISjY
GioZ6LVF1/h63BbGerTDSTQfOGG1JyP8M/bbzolUGQn8jhpqm6JvYFnonbWgFo2xGpYSSuE7QFUQ
dDldUMwGrx7F9/QYJRJ9+UWpIk8IWp0XF4xihA02scuvaBlmuxKYlQyuVhPg/GRq/Dl9Zg+fAMSA
1Jsflwt7ZzQtY3zAa+BcbvrnYqroc0sQQZgDCBj+IfAXw2FoIKo1DUMcVsCjMoCaIt9/DGwEN+kj
HEuOOeN4S4RzilPglk4b2R2h/uqnX5pwalqhgUQPvbUHdn4xs9rf/SNAFB30Ue5+2M0mxwr2zDVm
xbRRKHYlNmyFkPIPIYmrhf2xOpRRDu249D+tbyPPPBMXP1KPj5yskli1zAtOXfSeadDAsjQkH7Hd
oBG4yF0i9LWtmwy4kL+oWex054hs7gPmUZ92E3sEY0CreadrR1TbYEy3RGmq2P6ABlxItTsrp6nH
Iv9MU5WzDcUyJNZg3GN7parhqd/WaE5ujkPD8Pw4IfYU4Q3n2rvCwA4oETufdWF2VPu/0h4B4PKk
yKow4up1E0kKqx7/0fnvKjBPv4RpyaB8IgQq7RMeBfd88cKQLSrdDssHVK3rbeYBmWY5gvlCG0ie
TQKCenZRIZgJu1It5yG/+cCeGf/iYA6OzqnYyJy2cPWia6K6IY38MWsH1o01UvXpXouryguN1yuV
HMSMRIkKygYJwjYQpgdxMunkl/5kDTCmGtTBvlTzjhBFcyPeJgImTd8idHIIw58rQuBXv2TX6X6r
QxmdJQse/cvzAbW/oDSI5T0QZnsCRoV7D6GMzSh6wxEy6cmUL1gLXZVbyzXuD9PEylK4lyhAVlNV
GP+SN3E3+Z0rYjuQm0zARoBuovkKEO5HvpX5gi3w3zaLZytU6P5cgT9Phut5onlP/onueL9wjzSN
PLLq1fYtcgLFcIDGkfHjdcQhvAJxm/TdlAvZUSS8NZoSSCOXCzqIsVncTApiUWgCi3h5BfCTXIUR
gY03xKu6auJeT/QCFhBzK5mY9N21nQ8OgTt37+w3iXKbFuWT/DOrgKfyDUoqsKrJUAeN/SsJ6oq4
lQGCkrWEwApsxhiTvQPIwYVcvif1CeEQm1KLOsK3VPi/hX7ptjpT0cuGqqJ/ehLJXgpU4CqeSh0x
+VdjABVyjPxi3hSiPRh1xx7zkUGeuqQdcIMcjZS73SvBQBrEYwKS2QemATmeT+NYmSWqCsYVC/vo
+RQ/OQ08ceYPhP5w66EK17neJ3tJq+2GhIZ8WmSJLultjmg0jM0blPQpa0aJIfQJQ3an+t6velI4
0FJYq8dz2tGOD1mYokjN3j4qbs2UscAHsfOhLiEFsR5EY3lbCssGepkuS2j/2ItkOONIx0FqFoSH
4LIf9Ouo21T+G8lDEy+M1jWz0xC0lwHBsxjCkW5yGloihf/ARr0/iK+UPHaBbwkKvtyzY9Kn0ne1
ph9wd1vMwNEOeuWV0gfV3eNUwL9jXBqKLQQVnogO1tiYcTeTFazAEVuxFdXQaZPNoBdkYV3HdeNx
2/MclZ/bdvHmD1komQLGzDrQyraiqaqC0f5y8KcPcducuRzRw3EHzP9ZcKZNrIzFuFwUM8ZhdQ/A
xX8UaRPvSQNmH8aRCHGD7V5WQ1SwQh5LH9CWvNO4FYkAzO++251BjtvQU+4e8KTZSJaFGYtbT6hq
OyqvGNP//+V961ZK+yq63JrO67WdHfa/KxdeoXEaY7kqiXnOEfiJtsoCkcpe58gGfiBO4UjT4Lyi
I6NfyqhKeRPY9qYYuVHRSQxSgYnvK45mk4wtQzMRPJPlmR6mPBM1zzDP6fdM83Hvur4mzOvaQMzt
X4SztZESjp++HTi/nqPDMuJcDA6ijpGsJmrLPUceFvB6R+5IFsxNqaFRqksmSon1HpbMM0ukKlBy
9guSo0LUaLIB6BAG1otZk8SaPydbct42wPop14GoBDOOc94VaOHaFgPWx6YORZsfzK85ZSKH5RGb
bsKCJKLhli6bRKdRJVY0cfFqts/oH/mdYS/wKonm1UdH3QNY/91iFVC21f9a7MLHWzhx/psHwzaw
f1aUKF9jL3S3YPRraFZoX7v2RqmSUlJl4oU2y5FBzH4zPGR9ygVwcV9tQPOvWHZ/KE3rgGRQ6JxT
p7t3ICJ5JU+g8qxxWcbxIdUailODBgsqWT2sNONy/SBgXkpN4hFt9jH6atKPzfxwSJMlLhdTwSw1
r0xsfGudI2ah7JlW/ju3Qqj6WMwe62K98EDilrT2jP1kPn97ZI1XLlpxs3HlBSoz5OW6a83yy5eh
NJ25KvjmXNCPvM0nUMdlEmcX9OU8iZuxaHo7/0WSPRuIsWOYpY2HWR8uO6M0nA4hc5JPEe1Te4WG
1XKj4OP00r6n7T8U7NrzyC5plvAPqrsp04g307MzZonmDBCBT6gP6z2zM0nxqczOGsaUMkNWCX9H
Lnyk9NtavLV7izULS2JlTy0p1k335Ii7AXFMWpYHNc9/y6xUgG18UFR2eAwrd/SfFqItX3j7FPoA
gM9YOqfEH3dwWsq9rtXnnW7Ti205kyNuLYuFFcDgw8ORyYUR7+dZi4ag7C/H+NLrT2ThRaTk6ZQK
NifSFqygxQ0oHwJ2KnVu7SxibHOc8mlb92bZw7as1CBTuv/KAkCkTgw0e/JuyQ+yK1IF2edY5MU0
H1ueqbIGCNg3okR/QC4a5Gaypu8dOm5Xpt6MhaGtQY3bA+22Xpm9BWGYUwlaZguhblhGduf4y/Ba
pk6L8Ybc6/6D9GGAA5e6UFsieSW8nmN48Ij+4toHY7YnYVB1L2jhrvLLuvmjz9o/qOpL5tHA7bWe
gemQtZL4QXHTcyRjf+U3Osb1nZvWm7s7S6Pc4RcdhKGvXzGRLW20wTlFoMeeMcPezLlzS14vIRh9
gvxI0bB+482uRFAesfXgfeS/e5QGzqbHr1I1CMalBawfNmaT6APqtLtdd9z9usuhYXoUHLds3s2L
zPghkpZRDALKWJHDglU6/0PYisFg/c4RU5bjIik1ggM17u7I0HtrcWc7JxwfqGeA6yDwwE6vEKQe
CsimUnYLdIFMkqM5Z5LVY8Lm8grygZptdteIOXYxjQjqrPhtxTebwOJTcq5Q3sMpAcr1iT1SKKXA
fI5NFY2hLJNyEGQBNiipWzobplO8zeYx3SiJIFwPXaBz/NR7Wl3KKLR+qUcUCEI+awI8ivivi9ce
hwmkNwPRFYnzkeaa+EBxRgI2rUV/kid65G0EZxuYwSbKTgMnnwIA3sZ8gLy5bgRcHnzDrfG8Jepc
c5xLJHbiBN5UfmK43qTMNIYIJ876md1+dc7DRt/7jPzVYRHagtJMBiphGwy9E3MRq5x0drqsT8QD
8Wk1rOzIsNP2qNBqSGfO1KrQ1kj1MRhxjqaJRGzXsk4uzmgdEcGZuGTGY8nDb8zOiS3XY4c7B8TY
AKhKSg3Svhf4yxIerIFvwEGXeHP13fS1tCOLC5WloTFpzrP/jA8JcX/5qDxfheAGIhd9wmsD4HgK
BnEMyZOCkfveyeyN2P4sYn1Q2PsCE3VJeS+bsoxUZGvhd5MPYX8Kp6Is8utLRQmLbHZb3nVGWeKx
BOem8bsLa/GiS2w8uIKyufE9Umq+dHdMDo9v9DVZAXn76U332Ot7Xyr5dALr+ytzRucCLz8BYMUU
7PyeuOguvAPj/EDgq4CH/QDcjyCBND7jB37VJyI3nKhzO+ObSaUI7rKlIUUvU8yHluEIKP00geeg
WMnD/DYB4D68nSLyVWCo60iA02IX3H5QtPs3B12NwTF0s8SGbo/d9NRZ/BSsTIxxYRhYbD881Jmf
8UOjCc9VEPMBNXqOLmh64BlLEyCooBYeLEIcp0FugOoQSfn++rogHxXbq4A6dICamqgH2zgEbQsF
/CIJ94rGxaFpxJuiWk9OTkCP1qKW4o/yeCrNNUq2O2eJe3YsCVgnsJLiWuJStG/+1dj/djnNwgk4
wlJ3BfAvHVT/Hc+A46IHsVlhE3qXn4holpAEFs1i9xIUht/AcUx3dc9LGg9tEymdeAiD56c+fxEZ
GswMzg/4emrSp+So6i8AquJ4bv+9/ykBXV6mqsl9nVRv6feV8DfyxeSSUQeFiNXFmgqiGRTyzaXH
gPoBboXglgOco6M01XKnF0dAYgyMD4pQoWqRJb2n8Uo4WDvl59MZL2GhPoESMBdkszfxXChbvWSO
Bifkcfr9nBh0tz8lvfwH5wDyo+w1Yb1DwMiRExhei1aWXMmU+FTZGz3o5h1ZtaKUly2vD7/sgxaS
F+pWBubF3U5qHyOUxcmA8FPg0egkWkZWkaER9FynuDP2sQOPCKMwYdCXiCtVDdYleKZqM+jJNzzu
MkQaa3gYRnX4oyfswPq0lQPtKXMR34yH8DGCTBYpUTqZYZiu8Wu1qaR8wjXbS9+ylpHRQSvnCG17
TR9aNhuQrzk24BW8tI8hZ9yvhGkuYvNHK/4Dv2ldG03i4+LI0hdAQMLdkG5l1ao+90CVtJMH8CoO
d+3MGXSskH1CFUyGB8bm/wdNWgbitoTY2shsMBV67gWg4K9XSDP/uOKeBNh+/jrTgCTQPF0cOuzT
T1JDGZYO0YLgiyUvvTD+Qojogot1i6EA1agikjna2L9V54Ihh7AJH9/ajT7TK2ozrL1wDnq/koS6
eSODovYOWf+oBG5nFZrbQ8bWZE+bS0cX+nOJJmJP1K/Vr85+AbDmYW1bN662rWoWt6sKSJ+GccRU
Pee2U3XmNWSQgQ/hJD0qQzITXnmIXtKg1n0V7ww5uOAW/6P2SvfarHRlVGmPjGdCNFAD16b9E7/i
5wdQlPv66CnftFkklEaDXuKCU5rcCSHjC6ViLZeocxniDH5J2TUjQbvuO9TJJzJ8e/mecI8yYgal
InvGa0EFdYXS9ocBXle6pIOw+ipjfECdh2dZ2oJM95QDhVq2BO3uapXqgv7G4m9tpDPdEZ8SqCAA
Pj3ww0xI7UI+DXitHAFHzk0DpRcS6qAXu2a/mHzEYPAYZn6cc6AdyioQdx2iZrEx29SaMRkPjduD
ADm2cjwSRHSDWw5my4S84qg5nyafO4TlIb30ccPYL7Zk2XUK7Lxdf4X4e014ml2rCbtv1oZhyNzs
Aiy+ccibmKyC3yCKTjJSS3r+KQPtMctZLeWSsjUNT/zGoR1XkywNdLTdWgC0OUrsTv271yc2rKfD
aSSeEaow+dmOhIPhMrOSoUykp0Vcff1CDTgnWJuTFiFU7kv9q+BuJiJmeZZUUxtKd17+Gh1H+Jxl
pZV7CT+DLqxjjpZuXgfcVpRqxXJbF6M0Rzoc7V9wImZR4N7/WMBIVMjnGwr0RwUFeVM2rI72z/FG
OC2YtVBIsFfd4tk1gX3DWYjcW1SXFxHh8YrA313xWKzv+0Vt8/6kNQnnWOKp5dSQIjkJhyMtJpkJ
206jdX1ho6Pg6nzjuzWYeus2g2iQF8xyiHgV0YPTGr/ppr8Mg9CRPFUuTbXwnTLDovDdKSFwlYyp
NbUBew9lhcwmfsOG3/jPZRpQ0Hk30YtEJ8P8Thu2bhn9DWQkl2GYaRrg83on92No691ZNWkeHM6b
OuV1UZrBnpVly/EXES88U8j39ZVHA6jSyyF92w15uRkKAkv3yhcJ8etjwJAxojbbWIQlzh1z7ZvI
aPoQMh/d+10Ui4rSieHvzMjQWdDS6w3d6BzBUBkiMHDyMGkf82ul1byhFNsfr4f6nrlGl/g2fFWJ
y0wCEU0fAgLoAkJ9xv0a5p5DinKw7kqX0TgTxtB1yZdA7DWlALjBtiGX5LiPONTXVbe50vXIDJOb
vmcT/BbYy6d2yhzVwnYPB5W/5EDptylrltZXttKwZU1z7DCSHAsVLLM7eg9UAb9JNL0NldT+nofV
51tRE1teYGIic+mb0VOyjD+IyyFNQ51WGk/Rb+q3ZCb0uJ56IHrgudE/HayNqEeVO7l212naqgtc
BU2bX7bmz+8Eu6qBktJ3y2j7XAZ72+cpBzRakepGKUrBgnSX6b3RBkoICeXPfKHRQ4tANuuwn/0y
S3Q/dYnWNMNomYQPfjHE+2riQoKuZ9v8k9SpoBkXBUCuwta5NlZO5089hMJbVldNLDWDGINOTGWB
6lRSOIHJpzNqMwRqI3tkRfFxHsfkEPw1F0lvko99XlufLeUZOQ8F3EPDNiIXw5RbReScFGVmT+Ay
BFq64qZLI5EhbHVNNM21FtWr6dkufn/glTKyGa1Qq+cylZiCGYZ5QDR3SfekpP325n+LUNFE03aY
k1JPJGnYE72vOAmPHvuVuTPzjma5ZZQKdMkjGWXDcm6JoLDmPuHsN4xb7dzYLQ9R0O9w5eRL2uM5
k0WXoDkTLNvHd+DnDmZVopncoD3/kR4Up0DMSblRWa8GlcpQEDEEvvcvfHt+cv1SKp6SoiViZSCA
TpqOEuAeX5yf77inikBu8upHE/dk+Qarc3jxZJ5c5yzwcMXzK1Kno4EDsCLGtEUoZ0gkBav67Q3o
3KVCRSt8nfOQy9tSfs0NuhsG+I8fiMLcvc8G+yJGs9D1+1gfpG3F1sVajfV3i0Ekr9SEh+voPwjf
OYI8dHboGAQ8XBaLp9vPfO3/rk2s+fJNzvtq0orhvMrRdTn/NRzP6RQYo4MNe+vcmhXi/xRaGW2E
treTXMU/8w0HLjM8gqjSGrzHFKj4xOwpDoNpR44NGlAjfUSkQrC0qxseIeMLVXPnJZaELDKy0+h6
4gSTi3Fc2zzB5cCQp3ywWp37jj2HfO3WMsQi7V2Mn2LpUlowB3HPT8YfrfpBMo7qAE6FPpId6hZr
6WW5p1WQn6OQ+bXq8FmVrvDorV2XC4w4tB6d5DXQSYxskgSLuyfoIBwaNA3lPQ46KnFuVqWW1yLh
0+IAsx49YOKUlfPT00CEC7Tl/RJdAcDoJ2ZwqUIxwBriHBFMdR8l4zY6z3ml56V1jBtsigdZ0L2d
nBD4XIQX3ZviqNm515jfHLwagaHyt8fYG0iqtvNjMQGmuSak3aHjS1UYE6+xr839suheteUzbWjQ
Edz9Sev6YMRVKdYtDprPoKmkGeCSP3Locu1NCmTdvn4m2h/BOx0zS0iJxPJS0b3Vfw8cTSxpOTKS
i+z/BnZwgAInb7AXllxyEZUIB0/uQkLTrR4KiKX0CB7FOUjon1hGx9tlq4xfQrUBqniQw5On2oG3
fyrmm7fLQrbupXM8kEzFb87jGxeWaCyAWuyae7Bm3tOXpKc+gj3s6p9q9a8DnToP6TolVs+g1BBK
vY0D3KB0yqUYJKZtYYgZof/Vty0lbgTlsA+gJnq8Bhd3IB4N55o9BYMDOvg6wv/X+dXqDNU6RaV7
ctYzB7bkHK2fYA83Rs81rZ1tgbUzsnecQoz2m7QKKhVHCWR10BgG89BIkmiUDFcWq40SBMhg9acq
bRPc1oYppUx2eL8XUhXp74Urflq6+Y4uneS/EW5rVC/2SBpuN7Ik285Mx0/DFXEaNH4089CSkPWV
5jdlGKfkAuZEgU8tSpqd9uDrm/6Pl/xFMCHkXrAj5NLdVqpMlUFPm6nReDZNcd8+MLbFJNCKpX8R
ZdgefDqUBruBBAiA+2m/geoaYnYq3GQ8hcOy8c0ITaeGkBelxMaVr9GD+7j6RgYFQePeG75Ua+E0
Y9dLTVIcKqk4XmyBlXGfFVjype0qqUm7DfXFqfvtr7/WtGh1KkfVlZGzfTwJDXgQuEwtXs94cipk
kIpdo5t0NWf0Zet3KdO9SGyaJ0cvkOHKtvGBSwdWP3GkyDUbZDRHan7xqjtCmYzZ8byOl6xxg3W9
rIOWOHM7kWTIR6jZkRI90x5T4CUZgdLQdD1JXRJA8N2f5EoG1lQsboWc85bvf5zWIzxT8k99gFY5
1dzutWIe7+gJ/YOaZSB0g8vFV1eFChzUlYToeC3y0jLX6XAnAdUCCSwIiVqJk5KiJ0tBIeZi2c5t
tDB4dneCZmD4RnMxbW9svKv2jYlTfj42/s/YXK3BGGNF+f5OksEgvJ3xUApWi4wDFpHK4vWokExh
jZBVpysdLxC+rvAlgRt7hANugtihBf9RbeZzxMJAZsORhn+tZ1SAKf9BGuivSqNbzfX/bni3gpei
uioG1UZTlZgjSRHrdUusO+LubP+NxO+vfKiFF793XhwbacW4zjUfXudYJ0OhNRqL987SJ4gbpEq6
lhfTo7YyXzz/9bNuiPf0jFcc8xbQVy8eLVVUPbHALXlYs4q/ZMzzQ96qaJypkJQyky7WMjK0lko6
Pp4IbZcppETFs9b9RHryhn7cQUiQWJnD5LyRZOkM1+8Cwv/U/scyWt20j7WXajvoZZx+VtRJ4lGN
4s/TJrwbQt0Hp1Xt/ozSFcHRsaSpQNh4vhlwRLHNKcGvBVcDgqBjYkhGKK7SJrUrLcGG/nB84Nrw
+DidwV7d+NCI6Km1II1BLb6CncuUWajRDdXjqnAv63lm8nbG3upw9rnIpsTH7QjSifwt2H+D94ed
BWGBb8tCLaHjBapCtWueqNPi+QCTmo66SjNJtswLb8KLsZBOL9j3lsQt0wQty1yppzmV4iXQzbIM
Iq0zICvCipeNZWwWCe626+qhKe7n1YHMcIi789c+AxeHcOd5VYcqQ1jlM/Jnh6+VXomOpIdSV+18
gc8KPED7t1EFVVrMKGUtQcWB9l3nomzeZi+zxVjjiBE6MSM7h7MNum34tz49M4Fx44kt9Wxl3q2i
ju7y5OvZDo7ooo1Mg/o5DiLEWCq7Rnr6I+QYQ6/GL/vc/VWi4x88W/MNQMjQrRDbmMN41dz0qT0L
STHRazkwi5Fvnqy6rOxsivjO2SGMOhsOultuz9AjeA0aQeN6hTofM0j2fq5xbsNQ5xOZYxNrogc+
b5OBRNq1sy7wANIrpdjuOe3faU/vMy64em98clrwrz7CZb7pOLq9VbCjsY07oze/ehcZe/8z82P8
bp6AKH8bx5wYTHj7kDqHkCpupNPEQmAILO8WttMN7JBdRLAGnQT0uC8sH52qGsbIiRww9VvgzzXq
JO0o1K+zF1ERkCqi86akUU5phqImV+kFVbIpGtDRC3buXRpf27wRkyhgLkXFe3n5Fd4E108Jt8Dn
ieEUBruKX4+LYd78jFqrKq4jBl9xzmbXpEqkAOeBEyuHzCekqqRN92x9yPYx2TdsSz1Uzetz83U+
PYbLlZDe9HiuYmTiRYn8MXTVL3nM6ejVsNd/ucXrylJpzUzGqRRBQeAbWztKJMDKU91mRJobJRxr
4rnjf5x+XiZ2VMSwq5dDdHoz0iva612G9DOCPo2mkgToNKdZ/BziQTOlD1yAJyoocXIZpAictlD2
43gYQMqFPvR3AZfNg0DiJoFVy+bJPo9SS6lzBD/aPQqEQUrjlEYBp31mGPJPPlqVY/Yr8NdpAtkz
IfnJ3Q9NZFEv4DM0flyKqILCaV9MZe4cE8ob+VLKtuX5yhDN9WvOmlexQ07jZzuFylXd+sE4Rwv2
v7nNrY7aEf5eUk2esdQih7YV03y1NkGMaSgSUhxZNJPMJXC+3bTj47Vp+rtJS1pI2V1SM37RoHHa
rh2U0ILYjzR7eqTWA4CJbzsPgewpi+p0+RLLHU8tBqnByKQVxHDUV1SZ3rEhkXVkVrtg4wu+WCBk
j/cvvppQF9R2LvL0uqVtE9CotQZJTLmQyWGpL266Rz8GoF/HdkO1hDi2WipVHJVtdbEYyYxEh36Z
6gQ9b2azICaMUEuGj55FwAwD9A0gmeEnxlChIwjgqlGNbcTn50mMsc4OuFa9F5S6vaa3R9bdc9Ku
lojHNgLjRbsMMYAv7YMX8LmwVrkqkkrfXswY/dhZ8jdTGx3aeg+SHd9X2oJmqQYg+4IAQM029xZH
K9AbZoUAfRpmdQSyqC6GzMnCHtoSEl2l+lRm37qwIwXuST93QmS/Ieow3OwTcP3MhCT7/eKxTeCx
TvVirBsn9ov2LZkEW/3WLNvNLSgXLxy0AcdrdyumUCaR49eH+alnXGXipJRigDNzGU97Q5AsgGku
Ca+f0n14TSe0Lwqbg5n84sWFTF5qyPXP0vW9wnPTFmawPfQudVIL28C0K4s35LVor4s85aumDrMP
aO9plhfxZpTW7OkOBLkWMNaOhbCUrRFiarxkdsLFvf681WkWfRh4I0L/YE3QarIJsFmZDMo37o4u
Ng/YsnWd8cvd5Zap9AaKI/DjgzTvGKnOjllVL6PV0sT/9I3iVm7jHaf/gMVTpbJatF2rIt7xJYsS
sSHXkcUUWNs4RyMMAt59xKfrKdg8Pd93y+n89WXjOvuZhoXG797i8x0EtaZoC4EIIGWQbREoJ+iB
p1fHD0qawjT0MIWF51JaPXEuX8LBmKgp5Buk/SqwOg3NRRTFbWVPB5XMwxkg253Bsa+n1NfOND1l
murjDGZuD/4suU4t+1Jd6G26GmoDypxvXSUpzXwre5dsodQbKWvzHjv+GhcISaVjBLlmygcHYciK
08lXYosi3q24fWPFHlPRpMGackUPfQ9ZyFLeS5Yz6CamKOjxDVjeV4qhXF4/cu+umlzqLVgTUql/
1CDLqN3PoBfin7XNgtNPbcEGmkeRUJF2e/ofoNIFEzVjwOR5UHWqyEBygb7OXrF1/9+aCtq/l7sH
SXNZZHz4hwt3b1IP17EiiJtlJBlmjjWSm+immtZCPWTnPVEBYA8K5sXiQHHcTZYBXg/caaJp3QHR
QQqZtI++icZhcfpZRon3gsRPihUnaHKb/G7ftFhjRWA+lrWjaRxkGTDSyr6ZPu9d/sk39R7xAriS
ectJdFbfxtuTGzVduULj44BTcPksAgCvRlJ6Iph9jaFpvkMYnX8QQPbZU8a7v6GZXr9zt5kRLgYo
dNc+W1rq45X5l/JEAGQXNe5H2mJRS93O52yvP1fYtwtXHYLDFHtZDGsRmFVGsx6Qd4ioSoz+SjLU
+LUo7BhzdYH4LgUBpkaSTPkKQUaathi13NStdYvz9l87cXKBuRp0aQUVTpt4Dno/JpeVAU0V0GwA
XP1fsyx8nRcNTWSYaV3OrewrT+eUhiVBrkTiZ3Jxz/o60J0vqi2qmwnelGDwkBSlABHTT4daMIXS
ndFpTsUwP5MBTV9l9PMr3fA2yJ6/a+5mldgCBSwPJKVT20B944BuHXxMJ+7vGZIQLDJgEC7/NMcs
w2p9u1z9w2urFsrdGE5fiGUezbjNHPibZQKJ3nIL7t7Of6kRB9TSRSrckmBmeZ4KHtIjI6GJkqZp
OCoVBdUEsev617IqJo76ZSPJQY6RadfoFzff4uxZw1lMGHrS9NBcb1hZxE7th7m9tRfVGjpWXAuM
r3cyq0sTf452QWE3rHdceY0ZBatVe9N6RuReXUjjneXZLz0fqIBip3QdExIa/RZqh5K5pTocPxvN
jDA8+NkrlfdcBLH2EN9P3ZpNjj8kXVAEQq3HLk2VxAQm0uq956jK0c+XOtSJhb1d8cusdhDKL1sH
AKSAfTJayCLRFkrcNtfVFJIMiR34Bl53OOziIOk0HW8j+o55xmsMa6CDPhZF5G//qof8ykEQmdYE
FMeZDbNrcjb7dZUIAXFKEZzZA+ca0GQbcM+vWYyxhih1lbIdvKjzcxfX4xbMSGic7iESKE9a5Q0i
EV98/RF1yptlec1kjivHajsJ6Sr/dlQOT11SxOJrNGTiWutdTBtFiJH6vx4JPQ+ZKOTIi5d50N/N
qNCFP2kExLbWQOzb9u4XWYxFAfHPuf3hDQ352IFo/nUFosAbNMbo07qm563e6EM2ItH8o35bL6yR
9Ai50+y7p9KK43xH5wpdBRM8pNlLemVTCzuyPYb8qKXpXPxPEUTLqDqurm/2PzYnHbi7bweWW3gb
AKkDmzAyXFNOz4+GbfdxlHwUR1v6qaLY/XcsrvbJRWzEmHzYV3Ec+feIUuh0JHJWp0vshcHwJKI2
pk181p12z33mAf+zQkINaPSJJ77Ywb8nNUFv1yNSHRVcH+5n/bRprH2MLjhU/o1n1C8dul4UaNgz
RyW3NAXMBnaKnkxnoUVmuKGTcw+O2ROTv9maO+wm04D8uoZ0dT3EQPt73Eco/md9ZG1sTBqKt1z5
tZ5HpQ0YG7BsI6g1ZJeh7GOaKO+U1FhK1qj7BjCYtLrkN3Ooq30c/Lo13V7ocX7o0apLWsI8Ig2q
DjucxmM/u5olzttbP4vjpPKp8Z7VW1e3/RRB4A6SKymc3M/lNnlfCCNZ6UQJsFE/P4ejwJJyzAnB
I4oLPDXDrJ1GFcxmMui8QQfRLse6F/s/p9qNblC37lIvDaNYZP8at6cLzabM6J9A+hDi/nzoK2x8
No4M8hLaP9tTXYVKVdp65uprUBfxwNhBjBtrq+bS5tmMX4Y3EuLq6zzQ+FNfqMNb+1iUgAeF8lsr
dOQWidOaZiXFMgQDJJk+PIlcnfHsXQOR1Lz/h1P4CNLrTKoRdUgDuBkfKVQ84H8dZ8X9BdmyaO/Z
cm0KDrzT7CtqHEMh0cR9k972+TlPhAOqBZmxHJLvytkrhCUyqJp2tkLNUy7xr+3jp7SiTSSXIklv
syAxvSf5owgdThn3/6FCffO3b7izUyGFIRmcNVmJmIuiHM3OblfmYuGk847KICUxJ5y4F996iuQG
LMQE6llmosAh4GgbTqcwB5BwnDVA9f3KzOjOHWl/SFCiY+Hh5bkJ4AjIz28RmlWeoc1fYsUJwwnv
NKHJn0fpFVpC9vvcZW0cA59QDLJMcDs39jO2J/KJsMdZD+Nj+8SfePah5+2lwixV0N63MvlSpmf5
ZJtYLuKr80xN1kXlUWrk3vYux5JsaJcszQMWCtsAPKCVo248fuAyx9hbsq7lmrOYPU9Fxmps0UEg
6Ni2u0ipvfHINo5NYh+TSYJLiNBL2wDonnFwhfslchc70Mz1yTfeF487e88iEYvYRVl4/ek2E6Xl
lP0JM7JMfxAqR5u0RqxuUGauvaee5VA4++64P+RPksC7Iq/Rk0M70osHtl9hWEGzUtr2NG1T2YCC
fCiyfnMPsjAQKjCD5traUKnRQMg/S1dqFOd4tdz+P0iZCOndQZDO2MKeSXCpN/xTJu/mEvOTlWm7
iT9U6ZjwYJMim8K8uzINqWUwbjNYwSyw7du+SHXU5CcCT1r8FdZV6DG2myiRyI+k9+V+GkDSaOlC
eByfeAwDAfd0L1k6RwHEs2Kq19g0TKUxy0O1iHRYD1sZUok4lxYoB0HrZGrykUadEaAir9kEuJnQ
qLZwdoRKPrn5yAtGB1O+Ki+UNW5yZo4XUa4fms6dF/i5T2HSw6CcZ339Oj8FKiLjb2Z8GVPGrbgq
nkvmmsH+HLIHVT4a8EhL3JZFWVHeyg0FHoGh0D9JdLIVu1L7pYxEBP7QNTL6ZAjJ6SM6j2sXET7d
JGzbASmXeV+qp2TTGX5ac+yiAwN44YvE5Pdzb2goDFt4pidUD3pkDsymVKXvkO9Cw4fRgVwv53xR
7GMeL4QNFMEryyWotGXLHWCr0mo6xky3Nl71bLo8Srp7dbl0BYwGRW9BI4Vt6I/TaBaRo/DdnPyA
n+ikKr0DfOAfquNrO9AeM+ijxxBLF2H9cupUADBM0f6Y9DMnGmC+Ed2/NFF9ZT4j+0ivzr4m0d3J
kkH/VQ2SgL2qFu4p5DYXE+ZsW/8isB7DkCX4Wt1QCbo7ZkWWO+sBsFeRVDeL9vj2bQVKWXKCdk2N
jSY8t7C6qEf2XtBnL+MTOnzdkmvwhtLffw+BDCCiDvmhomUHElJRn3CoKBbMqsmrUxDDz8vGyVAv
taWUAd0JX9dcwxtUyQW7uthANtbHSQLFVwKz3Lavs8CPfXWBarBG/wqEzp+HwGmt+FYJQWGSg25W
rw2WO06zIzA8+n1iJEtpcVrJeDAnPq3DLUIQpb3DRXt9FvTUCpZk5vAPqwgsvRoh1EkfmUoMj8Gf
Jsppx6IeKBmUR5E2ek9b3RLhmPVxJr0COjbDZF36roD86ark5jrEh8yHerDpiCcWUlXSqr4lXVKD
/mlw2D84nN9hwndhiO9cYVKQmQlqETfxAGxgKr9VX2z6J58ezZcepU0vSSVsEeIqdclKIg8GPv1Q
lOyLa9lkWmySaX3ZT4NT0yv3Uc+59z7s6amGWqxQG+DuzVFZ/jhZ2iYVQF5GKvr4Ux0bXYQw4+Tb
b8hfdbhSz6MFmEMXMy5QBRwbimPUdEHu5rYNq5bMrGTvOA9Kp5Eyh+zYEahskE+cS8xMjLBAMQSN
DoUE0ZilRuzLddF4M1pTKJVGMwzps5kuiawM6CcQ7u91ti0186DUFEGQMBUExnOuKLxFxsU/SdxI
nXJQNFzRv/xVTPvuueUXNhOdMTKEDKM/dPErCLVlc6ut7XRU0re1vgy90srZ8/0IcU3qh2DNt9ca
sJ62y8R70Pd8xgisxcMwkJt/7deN5WHThERG2pMROrnBV2LoV7XofI9dYuA4FDwhjlmaPp2JVj4u
i3BdKzJ+XPTYvBwPjGVgkzUy5Uc0XSekBXaIQovGfGU1Asb1XlDOgywID3d2YNlcCYnAR7cqYwWB
HAGV80Hca9Mx7aDbJSDQBnrzFN5puPcarx1FIS0zz8qgW0l4UDROi5eC1FtrHLM9Ngn+ZJsV6Wjn
3aDFCxJuJNHaD2Q0Ce5nuhWnYluYGVs33srFl9jsXtBU6EcTVGrrq1smxmEvzbbbdt8/TP8e9nDG
ajDQbaJyI4MasiO0NCKqvzYupeF0CQcSdyMYFrcPBRc5lttD6zRY7Fs7QDYiE82iErqLpcr/eyld
5lwcxZBRsZHZoqGswquhCULnz2pxaq5O2dI7tTOxXYiG9Y89doGRwWvPYue6Pf/ulZAyJD1ZpnXA
SnjeiwPOYNi0zNYc5xUBfzzT2Of/qKwNjUncILkiGu1zv7pF6z2hW1XjnyOgDz9Df/I6kaL/tSQ/
nEAJa6klS80xnzAp+v9fM3Ti0to27yf6i2W7+4EY5ru3JPaFsOvKih2/jYaq+b3VGrD0zUJrxh99
AD99YH9ocJcgHS4GTtXC68t89AJd/D9RY1Vdv5gtRAF82e7ICmQ5yexZfbvZKnm31zpxBJMJeVyP
xiJbNye7WD8FsB2shnWbgMntWO5tQ2aHw2PgWtxAQI9zA2f0tyRmAChFcDdYFK4XtH5zBialR/eE
1ryfYcbVTcc/b8NueyQGhdB19UUpwe3I7rRndo23L7nbeVpgbhEqDBuAjXZ1g3JsddtGh75ev+JX
npuFK7efO/lRthASuJjdw2lQcA30XP0dAm0eMiyjPkuL8whdBzRUng3SXIqm/I5fniz3mGCy+wtf
R7/JznBFligTb5YRIZz0z6RvJ40aDBFXv7vhE3XNE8kuTf0MLaV3GpA759WO8VykXJ7TLfubv/wa
TQFdIBVSbYhxYBMxbH+dLhH+8zdPJeb/L4KRlDN7ZNUYHd3Jtp45Br5QS2roZVZx+w+rJDYmLv68
BbCLPDYUJM7LdgRjVrhWUUgYtnS4r1JhLk+As4Jz8igbj29ahcG8emjYKdgeza1Vt31gk3cJGGUk
kKOadpcWJiLcpZ1j1hWLr7JRt8zs6hWM3GwB1T1hbDMtRpIyIcLRZmahtCNUeYBeLz5Dwjy433AP
Ch4ot88j4ICKvYKN1rqZOUCGlXvQ2PVKp3nFWhEykauVMQD8Y4E2Ex46ZLBGIg2FRr1fssNPg36t
ipx60oZ02dwPqOTABJGNRf3QmGFJtkLszfgI4ZWBR9aqWSqpEV7ppmWKDWXHZ2jVQDPrWII8c0tU
x0o6V04f4XB8lX0yqeHiOhvyTcRktfzVZmwXkFYqGQ0XKukvzVzJEdnhAUj4SgfZB+ZxQVSIwLeB
wcwXJnN0ggSePm3kCzlvm1NmrZYGd1Muj/hMyQLGtZ3uw1qyBt6zalj32BPy2NyByJLH/1qaVpzp
7SC7TaIhy/Wr1n8L3dhHaV6UttD2bwAazy3Kx6JD3kbsbBvr3tat8qbweQsTfsqKC8PH/MSIKw2d
4Roqx1DZfiq4zyEux7LgX6rNZkVIRmImpkoDxo4SQifHdWR3dPqsQizuGoop+hWVstgAxjfSsNXe
FZ+prxG+3saUe/Qlas4a8siJVja7IijRsKgbdBhKymaFHCBRHFoSkZ7ljQXQ/acZRbww3AYE5Gu3
URcTH/IrJTFM5vssbikHKTeAGU1463RgT5/2kxpaVkGfWFMK5iZilG5oz3OLbUu44ei8Lc1CbKIU
qefwGYgWSvHTB2ZDgsExQ256FArrceS4KCI7jtZRNBcCHNgAE3JdJwOcGrlnpupSpRJWOUFiz5xy
zc7LG5/d9PHcn9RAdlKE1H/RQ0Tog5Qso4IDCgoi/9GJo8SF7eTr924DgZ4LeVQVRGdP9aTBet1A
1RYUYQ1npYxPFLzWCvTkhEfWN7jGou0tIu5X/ivZPYVHzsc26aEzR2Q0EgwMTNg+53MseAnYX/Wt
NzzJ92IJUll9W+4waw4bGCSHFDlx2qJsQq0LwmJgEmlx1vbv2j3sGJWguWw/mH2+RbByn4utXKgl
A/FjWx4pkURyKbLIyX8FmGtawV9qBaUlvRU3LdmHX/R8/b2ZKLCIak+v8rZ3hde1HKDSbUgCPdgZ
I1WzCHOXsvq0SOZuk2b+ldUXhlMVdEDqpzdawK6ey72Q+TadlpGf8/oK9l1MK11m0I3olevTRQ/O
opEwzospaTFmElZCCLmSCZ/PSNrLrpj3b8OhpGCW/OPwvXSUVwdxUgkRoaZ2itSCrlwnUkDbmkCG
Rv4oHV6Nzjm+EXI9RtYHiGlwHoamONgdIM7ySSvs15pQO7Mzgthz2ZBmiMYgyuCG2wOHiLDG8SOY
t/OQhfoxi5mu2Dmc9QZAl3kmVmFYR8L0qHzRwPbzS/34XR+1uJ28PHtLpZFMoFXtJ/yQl5vIjNhR
b1cFtCZNt2uuNIBx1I3aTOuRjIkIslWNZByDoU5vP8mkB9Iu4Upb1fc3EIcaBjj/qfZT+ME6UgDn
HMyLRcqHdaylBxMz+c1B/Fir/btCWbtNm/2dvDXSM7qRvMjJQZ1AL7Y+hWyf6D4WI/aH/EiLWUZX
SYB61VjNUZizgN3mFdYXaZF4TudU/ZYydLL02jx0K0u2WuIgo7Ij3SClRXONUnYElv3ebAVYutJ6
sW2rjZOUVdJD0A3i/8K/mkgi0yM+X7l44wEuAUKhLn8L4u5HxxLeSO5w91gLZdiCqrfE8ZI0RKCi
ll/S+v1Guf73vWgk1Zr02PYWGKxt2QC6lJPVBlSu4z3teUJrMue1qmJZWBJ9tpZPerbl+ANBA9yW
62KYT3qk+65LlS/OtO5n+vo0x3+PzUZlw/eeajvLc5wWEeBHhfiMWrkgfPwKCwcgdEZkG6D+TrEE
0GqWkE+kIT8IBTphQ/vO1sNIIi0ft0CaSGJou4DeOtp/QWF5jXf3hSAOY5XhrAvUyBePLkE9KQnB
L8GUv6RIAuDn28CwplWFWhxZxiKgQTyN03TXcFdZ+iXtS9coYBwpADGQqG0vcYujatEyaDbiLXbL
1mYX4KKLFLsDRnajR0AoVDXnPvs353hBmSPxgK3BWNi/GJpR852PumQRk1SzmMXZYTyEB1TiV92e
ZeeKc0Qm3r2gZyRYfJw3ko45i1hlXBLuORzM7kdFkOqveUahiw8rSbB80xbUALpfqNTx40G7UyD6
Kj9iuV6uTCUt7CZ+ImflsyyC5Pi9gUvMPDk+zmX44QOfi4FRuRnbO5XN7dWKpPFzWaT7yoqUoTh9
GPD/5n1CLJvWZEj7o1ii33xTkDrp68vGMU47dInPN9+uQwcIzXKnVwsFA/+3Qpq1b+e+cb72FwAl
AjvmFUTesvMSF+M3CXNmdFXKvpoXI9HSCOBN6WYtAETCHBxrWF6w64aFI8Ted8YggE950ET6yoVd
Z4Csx9NaV24ga7goLbgigj7cVP4AxLc/yFDSyE5IgFuyUzMvVH0Y00br6gQwXEZKb78vpPGnDsyY
O0mScOscxzOqQ9CveO2ivpLcEgRLyoXL4z9S8O27NYt3WuCMpILImhC0YZWgERFwC2lBlPVqakbE
2GmRR7DTOCwwZvDUb/s0RU8xlxe87E65xstJCZnMgV3QJ1sCWgNnNLrfMghLvUVcXs72r0zLh44d
JMPOLpphmwCqxOt8WOm3qpnLggoGi1L9nP16FFFi3UFvfWPK7grtgE8pIq41LGZfIyw4rxIxY91V
ezd4LMpeuJ8WrWW9iER7FTsLC0vahZRUmuJiLeLAd/bKmq2Y+73bcXp9RmebjQFpq2/cjF27TiPp
82GxqvCpoOz29tCO6G84J/Oki+NlHo4NeX588EO9KJ1BZeAddQTGfKihUPjxDHTKPORf4D3hKGAS
fwDJyy42TGqEOR3KLoDN+izOpbkkyD/ZFdVE68323zqzR0NIZ1KOysByUPSUJ2HaVf475SCikhNb
uAZjS8+klMOGl0UnvRxyy4u0ILzqUv3U0uEA5q56neFjLhM6kArlwqO2VUc3uU7TFWEXZzysnWUX
gdOz2tYXB4nY9mrQeeT5yaJTeVI5Xby2DAhEsTn+EsRkRp8HDkjbhiQ/DLQlcxpDI2ILrYcfBpVy
bY3ysS/MXmo+prnrr0ZKeczjzxkGyp/t4NnQuylVqqL40uToRgLkVdFG8f/zVxni+ztsEdsJMRuS
Ms4085mS/nG70kmli8x2gYDE46ChcZcV6gaumwN1UMR/8cP9lDEHPg4hFZ147nRnOdaNmZDBA3Mp
bvHSVcNQjSTsdwmyJ/SILvpbwyT+0ww11Ufj73dkhwRXYMY4u4CJ3x06On1RWSffrtHasp8dXGXB
FUHzlhCqRMpHCjb96iF4oPnGJSLD4u9fqEqHXQE9qWjeOenJQBn4t4hZMnpyGuMKGgqSrGs0RImY
QWaPDGcYzUE1ecOGFOfXoVUWTSn/ZKQHV4goQAhNLMBPrLEZ0a9b/XSDRow/IISApTlIWHkq+Am6
Gl+ct3VgMDmxua5v3bMwsVWhT+SsAWek9rqh40kHWcSetwSCfR6BMX1Xv/P6O4PEcrrCyRnI3611
ixSeZvRn51UfZfW0m0ZIlO5NRoC/n9KS6GlZWujfFEfXgG+Mk78epLCdfaytbOYHtk+pFb973w2/
vxS0swz/dqX/8e6Yl1vrQQj5R2lmSfWPLfXXoY6/Occ7+Gt6y5UEFEhzKcKtC0CPOvJ+vbvllkq3
3OQ+Wv22IS4ju3YAXinHSXJF3cHtODjGGsbkChujtr7atpKpbqZfktxZcc4ZYoktrCouG6iSz1AS
GcIAVFjFjhCVbYKuURxPwoF4U1mAAjqHIM2mmundUqPsOIrRyesh0nyhnAWAT1Qfd87kxaRYj5Sf
h1FKZAiPsK7lW2cbrCcsG3y39PTZ/bIpBp9PqbdZ8KDxcrWuPXxbg8xxhmYYlBqbnFF9aZgl0aVm
BlbA2G//IOTVUKbAluPP53+zOOW9izHhfIoiOyG63eXvIW+UTkRh3guLRnxGjB6X0TYmk63FbfD1
4LAsgUYV1iWz/MsmLUT+VKsPthTFzcTikMzpnwavmKD3EHXhICWrcftzdz8nCVGhYHRuY6j/qvP9
pC7AN5KR3TOgHfl38E8VwVUrLPZ7uAaRqngXNm/Vf5kefti95WqfvvrXQjP/kQ65NfEfyLvLUNng
9BI8RKKmvImgXt54IC5WiQQwgrO6Srrn723EsXJGbL8AOPMz6UyxKxk0QWzZMJi4FnOAsIgkugZa
ePhg/cWqKeJU0FLs0GrMwi6/36dDt3Sns9yv43/6B3/H2i/9qO6b7ZJqI8TfswCdinNSM2fF3jGy
fDTNFPKvUEdctN83Xef3ohOkU87uHhSXEAxSxxfl5C+vdomGYQehxczv6DrUtyXvwM3aSBENL45m
1aln6m63SWLebhQ6gPhz8l9vxJiUdpcqwIBDF41ZdiI5/sXMMHl1nzd5n+Z2U6sydheA05Zq6Pgi
4AgpEOeC0XfRvWkA39DF4fx1hQtwGRg6A3nDGVH3d6TvnC/HV6gLsqOlv+ZzqiwLr0ZdForrbufl
VAgZG2NKLlfTwm8xqRcL3N0/1lGZ6C9aJudUMVP/pGwCGW/ayRPbnlQUkfCvduGxZ3iGzZcyhT1O
NXbz4sgDCbAN1EbtQB28uRL+In63Ka9AVZoTwfAjiVfNc8UVvQGPlJcleF6Y8dv8J34wUl0zt1H0
D8y02qHPT+t1eHO6x10bVI7vap7AZNCZPU7I/u//oZq0lwx9VvYK2tshTiw0USGVN9h14wilegqU
GgZKVxRW8pMrjeuAIU7mmRTjBAnjCHi2vP9uNm0z9L6DDILDdaePT42Y/ugNmeBlEnXodAf6WZH8
+ibKrLYJPCorBmDM4LeTXg3VjiW/TdAI/ZNdHb5qqCsQaG+QynMQuWKMvOIPTBXqrDYKF0f3OCb0
brbYwTofS3OP0kTzhrS3Qt7AnpmqdVDMR3IRex2c/VmO+dwxHRfpDWVcMSAcPJXIc545ZQPF4xK+
Rtz3v6phqbVa4/EQCGXucVG1PdgkCWkpdLRa+QnDaTW6MEvqE1hmcDwe0rChsQemcDy5g4lmdm3n
IdtNMQcGW6rqLBtYXTQACM6kB4lj1ayevqu1/OcdrkhrBe+6+0Nz7qJfiHm05ZdPwmRkHPH0hnLF
2SL563u4P8neFlupmrG8NXnTf8DZu08TpycwWt0+Sh7LTpXYlddDfy2pPDYL429lb9Zr79iRBhy6
Rpn4hrW+BCXPbAghCpCCLuCoiLtX2NQ7elf2Glfcj7Tsa2egLCwvtHGuS6EkmiMEqFisvrM207N1
NLHSXv87Uz8XaBYYu692Q3wVpbD3rPEmJZM3dYb4YTfeL2a3gPw4/sd+F4FQLbWDIqBPxkqNR4zr
D/YymM19LfMfQg2ESzf0RBG21tfsqcqLdMMErGylPAO8tFeaVhRPpF1aB7UGdFGRVfNz83VBXSIZ
GCabGgm+njZNUXorvNLVtUEuA81VaIYFZDDV/x93k365Z1yZy6LQX5g/ueOiBjPpHQzyzONKxWXZ
4XY9qXpgIHzUhAe7wbBLnQkTTTfvWMkiaCsZEjlDxsL8ekWAGp+9Ep9KRywFvuBrGNteaBGu5kNS
mxyKI+5VS2qB+FBar+jV2e2xk47UGakKqMLY/2aA1X2hACYGQNYbYvRkNDO5PVPgvtg82Red0Crm
SYDGGPCOC3ctGuR/Ye93ONemRFRFQbmkDFsDFneGZQGgQsyv6Dn4g2Kp9Q8sQmnSlsiL9tsHi0pv
3lHAheUn1eQzkpRXjkTe5E5PeJ67s+19KVQZmD3qtL/MyZrApz/nw8bYkXCWoKUtVKH7wFH0ABSY
D3go2an4cHhbTPXdHft3tMf3RNsvVZfJLgYWtfExb+xH2dNSQcsq3+A9sqhDnTzEAa5+uO/oylDt
N4gYxtgARc7x9uCY+T+HPCrdeZdR6MrAxsBbjuIBF8u/KOBPvXTOjo/sX+67FP6oYyk4HQvfqtQ0
Q7PgucQrTpLxgCkeoovsHDqFB1ATnvjyq2wC9/xOB3zgW1EX/cOcRENwBY5OrDneWVKM150uebJT
oDEioYIAmgC8R/6f+lMKG+FQuimdWilJ+kJ2Bn7cM7OJpNHrhAfcLzAKGYshhGbwiZCWsFpwHp91
spfVa4Aw4bBYUm4cT8munY5pjgXfbTalNw/wqz9bwpWWmCkpShDsqrrEMLQHCWOW3tWENC7kGxhy
tkgHSekf4bd2Hp4FnC9cvHTN2zLjavpUPaSu+73y4apH945UZziXFoIutktTFU2EigWr7KyPHwmR
ns7CVzi5fLotXeOHgoqxHOHpQLnZnpYE9OwBuE3kAoCoQnU6Gt7/8qKAxr7+chg2GWmnfPBV9kZj
M06o4XXyl0D44RsiFATbC7AaVVdOn5FgKieOLqrD+8/OwoEBmINOIyVE81zf5c2wAoEU2vuDjsRy
2A7gDTk7sZU2+WEUa2svq89nkGNmd3gGC9BSbBy+qggh5t5tYOmBsXbU6h5mIllWevloRNR5m8MQ
dhs/drMj+KVGMbUYZYiezGa+8TNxPqAmrqpS8qXW3De4nIOwhSa6bc5CqvgkRM0D2xzu/ZRXHjHQ
+Ql/NXaNHRMerIFPt5yJJqNkYNxvODszum3jjQPRqunLanH1NOeFcyNfreOEu/jci3yKQ9uoznXH
1BaYVxdwpmFDfozYGy+FCcuoY8tNPvJN5zKfV6AQl8CBfOyh1CC3K05QKMF8Pk5jl3R1p7jiFJX1
KZkvZ6CVfFw3Zv7qy0mIQr4TTGAVn1DGH7r5raxo7JZWEZSs8oKQfyIHouqKqdZEDNFfVsWG5RRF
rDbe5qL3NPcTqK48UAE4J3nGwht1JJbavI8MZBl75FaVymJydtCE5vT92O4CyQQwNpATw598sqfk
UCaVQfx8gbGIQOTmslx3lqSbn0ezRVZLvw9zPgkrHbzjWnY9uNFK4LmATsjWwTLj4miuLJu4mPou
D8CmeD4FJjTNBl9s5y2MA0kMtbqt1ATbn/gs0TjihFgqPiCjLs5ZRFg2H3K4fA2RD6W7ULdTq/gv
NpETjsJz/+WtPfveSih0cTeYbAp8skB5tnjusv9Khe+3sQB/sY8B1mCCTYT71QfwRDOTo5rSKQLp
DY75BNQVAKqwAbKsB3IDwzdoA4o4B2Q/xhRxdsH0vOOYVLnA7BaFrbqEqQIWIYwHkM3UFHIQavP8
ZiXu6gXle9gVE5OsXEcZ4LhSPYIgwPuf3ZTCpGkgeRh/wB8y2xUUsseyGGmaJSXS0BjQS9kYNjbL
RPB8pihkMI1ZbIZzuxQwatLSnd8XuRMa3EjZzEZMmNllWVPgfwzisknJ8w8YVRW4LuthyHQGdp7C
Oei+hLBCOprfLs71puZdzGHGEtTZ4L/xz4Jcs4Ww9J6aX8AzQ6Ua6cswSu9ugPIUJ7Hhi+rKc8tj
4A9OvpIS/NZTBQEQOwfOGBrtBJ8SnwEOAIB4JivJZZ9xTo3Eu1FCZJ2ndezoQLKPqpy4ZDXn5qIi
hMg+KpODOIIXhEINaC/Jat/SEvKPv7NTAYyfpbqwqw6XS6GPTb7Fmp/WHsZ0VGvPIFf9z+6Zam3v
smp8ndctGQ2OO7fgjQAvN7tFzkcullrrU38ltOYUCS59meOIP4T1czQgL5P0//mEPfLj2GpJlKOG
CMXl6USbZNuuyPEUqgRPOlkKU3I/QpPokMfDpy0VBIEHElR3JUApaHjeg6Jlnxg/B2WdST/sq70b
OKJqJZN0WTtJT7MRL6i2hXEqPxKZflIFHBLHA9gcwSctRhRGs5HF1ABqi6tzRf2WeZb/fXO8e9K9
RwNBgOYyrxMftEHb66uwGpzFiGXRS1mkiEskFdi1CzNgA2KYjY7MfFaLdIlRug+rbT7xzI6Cs+/U
E9qT2YGY8jPNXec3Fr9/ILqqZf5b8wIyNDOEIuDWOtTE94ocYGenBYOjr2ejAuM6KVvMWlElgZof
+l1INWaDfcg8I1BBtSgdIYl3aK6CfreNHMnjfPvi3AdQd4Iexp4K9kL0QrttMtQqX+8kYCNS7cUI
Ylj8yjuF9cMa1eVuar6+06rhF5U6aROUftLo/5ppOF2aVXrXnt4PkShjwDlqsHuORFdv+DL9s0gU
0lP+5rxB7kmxdtTCUTwAWDcpRMlCow47YOmliMNCQwNZWC/p8KuvXxnlrtvMybimtfHlqxFPOqVJ
+mNZ5b6DpEcjYMRfnzdk7YNCPNG69Q5zfv+ryBjKxyUUJJMl7XDm1IO4QD7BpRow8++FHoiXU1Oo
yS+yfQC/6eMPyVgIO5cyDsvyjmRpYBhP0eaofujF7ocaUh2yPq2jPSxtm9YLnJHiY9PwptI6PqWc
FTAyk6ikYApqzHIyYIRQoFDaFA4HJ5x705ygMgYvu8ok8be9RsZluNGb+HAtx7/DcSEoDPr9ynYz
wPKNkxrlOTYraaXNX/5e84DuyRc1SUHhl2QO+Ng6y6bPeSajqVk3wD7nh2DuHcNJTC+kRAI20b82
1V5er0pTQC3LU3PSD60P+4iIVrL9lb8XDH5FZrpVYX8L1NU78cBuUflr1pqajnpake6OHW6LBonw
ECvdOiwmtZ1Wx3BsRKvosFEd0ZAD/BrC8tS8fSRXVywwjAGq4qZS0QYO2zkpPB+XCn1ekSP/ClyI
L99G9bzj2xeLlESHi8ThEs4iINKkCHEKVrWYmJVzFEYdgF0PWGmQFsQEUftBN08KQjR5jVdr+o75
7Tha7ACyRvrmevFoIR1KRNZvFniLVML+nR4fW3qr5sclCkzdgmChUmBbGsoHg5ZckqjdSWWmJR7J
66vwyWeE9/4Y8kMaxHMLqe4o85ublK54qzcbPG/RkYantlXMKAsVNteuXSq8eQNyxmVo7icywrEU
NCMb8FKbtI+cCLiioWUjBfKbBF5Fk+CJgnM2hxswWj+sySZ14Ozl8Kt9GKyRz946YygcxM8lFAjn
FJPNx4UfY12C12K1X8iq7Jz7AOq5QkUuZVOfVqikYwxKitShWn8YssS3pTY8U9UJrHFUjh7d0HIC
IW8lTMsurvaBI/OleW8qhE1yar5W1qm7moLItCJRDoD1hGLbhwWTU3SPyDMSCysVrXBSny3EdOYK
3rfxBINHvgb+3H5z2osjbyxAuT1Lvv5TIq1EIMegOvNgwht70G+bS0LikMzir8wGstOMeURr/CTm
xrpYXx+Tjsoc7Q+7EUNt/phWX9GHN4I9KKrgdyMJavy4SKFxNWcGJbQYbfdAHnNgJTUnWuApg6gD
Z6tb97rdyreZs24o/gqZnAqqgIky6oyybzvVtR8WOrEh30D7EsK53Zqdl5+jcpnqI44rT71UykW+
smVOKdEtZ/mdqXMgDEKTnGmBfFaiVlIlWfvK4K/Kee4/FKe3fLOdBLWLYwWLRAFTs7ZwQGkIoloT
HAY9gGsrY3KfbSzETyNmAQNvQB6iNdZjScoNMi5Ba7wgV4FHARjYPDFit5i3zPBIuTU1xD2TCxHI
w1uzGSDMqkZ+QJSKc/yY6VFfHFjSF/f8hpjF3LAAtXJB5KG+q9tivB5Otq4GnShb9PYV8RRFo13+
U9ZHpb9iPu1Ha4wxJW5AkD62/K9t7MKRxRYq3dsaW5V1kUBOWFai7XCQFZvSk6dP8ZwtTbpkQb/3
zyzcI097T/c/dHC20XDJnl+V7II97KlBP4Pn5ECz+9QtoofMACxrW3GK385E30E8ds3Xmrhdg144
rTfKqoDDXcM3N+EveAB7SHCWObFnfmuAIHIfvdPdHkeYc8khfYQc9EsTOex0A+jbopB3IneJ8WrK
fWSLtvXHqJDRpErLsicVsqOOuYS5uwsdxzhcFjedLeMSkcSiOjnVx81UscyZ/GMjuF/5vwcdfyVQ
jBphdip6lGTO+HRfQFKn+N45J62O8S/ayITOgnnh648Kwb/Gi8ezUEn/KJpFRaezpc3veD8wnTH8
5z0pH7LywTsTFLDX7kqw1Ppv9heAs98ir1TlUqy+Wcl3ZUcNR3iLpuMBJz6VdPsTUZFx/cztcFst
qMKIRX7xL2ojiogWZBtym7X78WlIBb8X9sluFwf+IbjniTllMegNXGEt44AsdD/W9Uv1WG9bO2rw
ZZ9b/8Wnc4uIl5R0ZtgGEI8c4Wlyfd5pW3FSzEXV9lHkGT1EBwYPtBqTBwMySiA5C1TK+o0Ic/H/
3iymrGiQXXiFn4/ltNsJ/uHxdibbchq90N67YMw2CFmL64DhTPVxal5vTYtddiiWUG40swFF3ltI
QI93kRf8kW2EYoNK2z/C4OygW0BiiSYPWZHzA7jg4WjyCJVnU2fqFnI4uABMurFtUt82CsTS8TDj
OV9Bmxt+9znGTrLbiDeXQM4qoNMeLhmNS2+G51FvrnkGLP8Q0N85fxCKzk7kwi3NYUS6f5QSiV0f
hgjmbQJ016SPhzm+UNfLSX5eomHaqkPY2s0sLgQNpeMk2oP0ZJGSybIVQh2vN8QefekrkwRNfznz
NKxMYzLqZLOSdOcStEdu6vkFKiM/nLdxD9+/S+wTrjWadoh8z4+ZdedoqKYt4mYKBEAk0DbftkmG
Zq5ng87j5D5hv81C2qvTz9Yn5SfKbRa1/L166byH8L5cWfSLFPLCG1GymZ4ASwAvQZ/gELBUlNPz
M6yrJWtZvLf0O93D5TYjcERA1T+WiuCUyaIBhJi9Nmfs7No0g3yiJqbfVCpuuHIrdeQ8kAQKHc1m
jOBPmgciNDlHdhADrbEEanzJOtk/jSQFp6RCvgkpQaS6z7WsUYOPGJsRmpNz1qoLTmGP+HzN0rjw
mXhr8rfzBG0v8ZoiUkcKSQfhNuEuLWhYch/vtuwl4nGYPNIn7SIdgDBqZYebtQDfVpnwJndfGM83
+4TdXdS2afmDxfnWkgU+61UVinLU2R1CBJdpgmrSFhKuWGy8PD4zQFXnu0bjOpvTiouN0jNw3I5J
sYOjMYSMF7A8/UI12lprKrDceDVhQ0cH0ienTbe56GSAcGC9JH4/ZBX10I8Y2PMhjw9Ietx4MzMH
Y4E63P8+D/x2lsRkJ20KsBI5EaeapDTwLMmZsH5oWFeVzKqtXOmHfmBlXeY/fZaE3AXf4u4oiDK0
kFaYANArCz2pja0WsdPKIFHalktpVrETdQlNwVFHGAMP3D7TcybZRj+MELBvmlURczQr9Ug/OVls
A7sYbfigy7usXqdnK4XA358dSKgWXmnDq9sDfFPzH5hTdEdQyoUjxSBmg4muaMJ9A6J2eCE3I0oE
2w460dZ5gSv2TPjGozzajyzR9pTRlwyKLkWONa1KXzxlBL9Atqnm+136FJhhq6owIVIvDgeXujax
fVBmSuQmJORR+bADo1AZpghVLfez6wXo767/Excc/45rgrZDk0P0Qc1VuLsjMf8SpNtMURnQ6aJk
8KWrV/IdTDlbWxEl96L3jSv7cPnI9Cq8ibLOCf6WRYAsmxxGVQkeFxAyGledPm38iPhRBQMMtPJE
cM69pCbSDf83RJ3+qY7jiJadHc5FJmiCUH33pHX5Fi0mX+6LRT3+yWhrSAhBPYveWKmts27pSSAS
DsH5xdIzA+MIc96SRiaf7KeLNOjwFbMg66yaUlk1RwS6nT+cc16n6sK5PWj2CWEd4a1UyFTSP49K
rVp3VJhYVEqQ+CMpZnkDRHaEd5FVPY6fDOEPckuNuq5xThFDKvHsAGNWVhpBf8mZRm/EY2jhdU24
5zIAah0XmDGxykScgRBasQJZPVS9Rr2Fo//aUnnxuDZn5Tk2D8uqxjxFwmqTpH4YOBSsNmvOdGX8
uEkFlk5uiA4gQfFwHgH7noL8ZeEPjyjf85CU3+l32tqrydQkkE9UoDyVx8TuxHcTjrEzLSAc3/kt
aufa1kN/3OxRz67FBXV+25B6fMUsFeD8DPNpgPWuPCzMYFk05xwMy9QbhL9iee7KSkVP8nLfm70A
qgREEgbxCgSpafqKjdBGJ70sLw2AXUzx0mUTETaTTJAE/iL3CGPpvtAZLk3jxgNTGWZn6ACLZvot
OerdVcEnJ5J9vivNvfDVyLMlVYFJC6yxgzy3B17k+/2Odia08mmpTwEJHGOmFSAO9UfwotpIq0Uw
MSSLCrOe8r+BFl7g6ha4rAnAPsAinjIuIopGYS2Izxkkn9ki2o8PNDpxXG+hjbV248VNMF1IFqXO
kq41qwa6jBIHmzwKcpNhyN0oAwNsvwJA1RRkQwddxWTc2PCCCI73TNmXZeEroSho3477L2SKDGSn
ucMnMWk9onI5ORUOoE3hhyf/CLtKxrUR4AFI+vg8SJEkBvJsSrrJITapVlVCHsEFfVOtQEE6OKAu
s7qjRc+2e7U/g4GfUtURuqns3S9Wrcu7uapGcInrcQR9LpkqVjmeWVHQmcMRU1PWG8KyvAnILgdI
N92/BQyK7xaf5FU2cHGm8inneCqIzn3qSiwzwmYDTqZP4wAoYNZ0cFZqnvQt1ez5e7oKb90HjLOA
jBpl/ogzja7aE8DowcpPbASMHzJziTsvjXgCuyY928xB7yLKRo2P1orOY6jWfa7kI1lhtVeQVyYW
2qcnpSDmDLtt3hYYL4k7xhWsNiL4Bm9vxKjXI7qSdEmDCt9KC2enp7xJYMR+3qfZtYGMBeiRTv4J
fz4pKFTKrxxaJie5DE6t99i9r1t2xjtxAQWV1Be74jFcHXYS5t6+petaq2AyJhuPz48Xy2ITC3M5
njAoPnFPe/JS6v98lYnfsexITlga1z+OnYglilJXqZ2JJcr/BSwGKr9kebaXv+GzxblfZfxxS1Yd
B9o0pEG2sIoU/Tbq5rTOEN6BknUFEPVD1nAId3QW/+MMzR6O0CdiHNGIIqSEkyqsV3fFG+moWjRm
C4Yy0Jh2YkVu6KJGl+dcMWww94ThJXFluFWxN6nEl59A6IfZqBnhOzAdilEhhFCI4hHEe4f8jrpa
Z8PIE6WUS97TfcSj+7xi4oK8pBA9uXD78N8ZVU7QFTeOHLyp3WgxIBAVIj0uLxhy32vCxfg8we9l
GiQlkvxTSlS1kU3qeGBmB8AqHbnGJfBEcZmCoOajo8jAHSlidWUDMc3UaZUFTM1za8MFrZHxXf26
pGIPLtX35NfFVSf7E/Y8bpy8a1e3610ymu/7ax+K43jtHG6GgqckEcUPoIJ7meajPSsZzsVFaynG
gWwtcsNuoQ1D4WZIpIos5qzjGFB7C/E3pk+t0R/nQFz2wFillJkeJUaUpXMC4QbJ4M/xkOlY/Wl+
DcKBnE8f/8C1DeIiODRnU2OtqpKE056dnYAo1s1clTSW4vDeAj8RwZMFWG+d9ttQQop0EEihiaU+
e49HhywCbmp5t/RkmtYxiHtCQvKOqNF7WTQ+1DNmWBOSdv3UAAkHyR4qfU/BSPTlsOKHHQr1V4AH
vNn0BZSQwx4/1IPovTlCFT+P87OAo9zcuDZMq6oL3H6HazXRBt88LGNbCmpc7lbHtzY92JmZX5oe
TzUkJqy9rWtGmf5f98/T6xacBf26VazJcLxvdqG6egCRNKd/us2ZPXN8KRU8XSbL53MCKB5Xt5mO
Z5qtnE+ePpUUxbTNxF1xyFJBUVtw+7osk4Z3ELr0HqKsie6UU8lgGMeHVcruCzPHHMTfyetJxekv
4oEZvBZhobDZRkHCxepA60g1tKDOFXteZOzJgrV2nPzACt6jjGjwA4zmDdRsuwTETFnor3nnwqF1
Zyu8knfmQGXy619sLV/IotaUxcR7pKEg9GQsxNdEPvE0Ppposiv27/fBpSTOANZLPQrjMVUtuGnV
aOn2o3YljTs49xZX/llDwgWskM0anWztq0JXLgZ06W9LdkdRT8uw2pXzE/rVYgewEBuuu42zE8xa
z+r8C6WsFHX01d+mE0BsroNqTJJn9Tggz36619O4bF1PMkvfaMg8VJ5J8ca5oAerxGzlQs43YtUd
VT6uHDPuylTimXuDgmhsjsKBrCk4/W4Tb5EM24K9ExEJowZfn3D3uR4iomFefAcPomwAr7kwreej
jeeMbJ0LO1HXRpC8Axp7numKwUot1nLGfdXOO/HzRRN/FAz14OsrRIRN4KUA8qCDRb9+NM1v29GD
5wlvN/fJ3AMRVGeiB147/KJhYkngproGRpBUFp4/qPFMNU5uHceZqHxdTMkQcRc+qSBvmb9e+9cz
E1cjQm3/ro+ozVmUt4kZ55mbgHWr/kR0YzMNbH8OMH371P26xcoHYuvrWBTO9k1PVezfLcsa85O6
fT0XF+q5fx7tdDWINT0YH5a9YnLknJ9wUlFKGnxW54afMcV78JIi/pCIVGMGnkkG8mnJloyXSbM9
vsB8b8bsOc0mJ2lBmf1Z/VlGkvwXdBwL4gBWjtDdTK1fgLp8W+NNokEZrvV6NojNbBDVsll44PGM
3MOSjQlhEMG7CprztYcBY7lMgM1RY1otW88A8DNOH7pZsBgq7fZYxL4VNrF7PUquac9tnoDhHIWg
YGnTWMjCQE04ncs2+40tQUPPTa0YZqsI4A/jkiCA2uBn2iR98MCPdW4UZTfIm9usD3zRFoUOwuew
JBhHjswTe0f21Ycb6emPBqQYRo0LzdESkUCmkYiW5bH9Nzsc2Td/jxN3Nk30c+N7lrQj1mhynhQC
FnXd59v8PVum0j+k+erFidAIt4GOh/mUTWymXJW5+Kr81X+fEWKmqUc9gKQHgmJFpRH0k7T51Teo
fHNtTWwaJGZBweUWwwLzLP2JIwSKl3+ifXgoe1YdrfYS7LdzpOb/lzCrE1/0STDzOe8wnROPhvFY
UgyfZ1RWNcVv1JkQwnX+UJ4WI8FD6cTVupW5OqkBvxs6Gvh708JWfgZ/PXBaxi1Xzi5d74Rln/b1
BqbDB+BwJ/nj3a/5KkwgMvw7nmngECRHjEVB+VqqSlXVJS5WNz/7HxFYda7sRyNk/vXJZ8IH2ENz
opPKfdM7f+e9tFLx43FtR/9dANqZUZfsoMM+KWsDe60W/QmG844GY4fFaI5n0dv/x2CqOmkRUj3B
NCk+OWhF03rJ3xNGViJsdrip368rb1v6ONc6CMhlFpzWttU1MRg06Isk1tj9fvh5Oxbgn66eMYY6
HaBUdK/Vw86TevdqKNDsIZkl3v5YNC/Mh4fogWdtSlG1KuDDrL7yK9MlY6X4XKHn49NPJGTQ/bDb
JIQKGGZtyqDKxx8/M4KDj380LVqubtXKmlDG1TuLsluKhOWn6wIc35qpHCLEHwcQC1HwxWoBg52u
dYa8+p2VWPvBK4BO2A1uozMOtWKw+zxV3thWegnFfexhMlHiuhO7qoA7jzYo930ZUE1b9EL5gxPy
lAj/Jaf5+CQFgL9dx2XWmXWK2kCKPI/ecGrH5PEEoxz5Fgjsct74lwla5ZoKER6fOZXpGzvuOP9F
edXrNRD0UDi0bxm0+Y2CmJiE55VcX8BmSRadbAGu02lmWMjNrtWrOImQ07iWx+J++rBp72BlNOM2
iWLkAouFJduYOy4doyu7n0PIY0vQ8ZQNrihxqaq/1wzVhiXTgX2OrgZt31eJaf1WOxjvy/WHupiw
O8aVrBLqEk0DFCvFJOPeM4MFNLtcUEJXEeISigUGhABBuSOVmGrSPMo3ju/cJV0vgnGLMtgbxrN/
dAefHmuDgwgi5GbKW+0L68Meozde/vdLcmjb3RCtyD+rtryFnKBgABJLUtxe+Dm2UjMqbWriR/ka
NMi/ByUHmUch9VpkWNQn749DF30gzCPSbHS+dNC2z8YQTO/r1FpKbe/gYMqnHIGc4zvgKAY+/Sf/
U4HdTB1kPKEmruy/ZbECkb4En65eQMFFmV+ojXQkyDBmF/cm8gLTobzkFo792KT3Q+zch8XrilU6
my8A6rV7qUKt/D2/8TWAW4jqr/DCMbdnEjr3ClJ0vMakEfOUEm1BLiKIGd/U4qyZiYE4LEhttHV5
5KpG6jFPub9PVJtXYPLgvxkPGfzvGFGlXpxBAS0+x8yIsKTy4EDqlIF/eK/QuhHPcEvbbo8czbwy
WZvBT3ohM4mWtmzACOr9ebWhGIM78/CcfO5nuN441J/OMsIZbNLkTWdWEtoN7m4NKy1XySn19JCG
9AXAgswW4kGHCmU2T3gBxocwtvMAFMwX3fYlyisVtk1Manf/k/KNU5s2jcaBNc/+hpQNy1Qo3hx6
v4+AFhmI4FqEnrQArx1d1d/dHvTV3xWudu4EGJSZjAsQl5XSD/OQqsIOgpP/LMR2dW3A3ExQco7J
ZdXaj4LwDDU44jn+gCceIO/DJR0aiUx+z9JjxXns/TomROuvrboEqhltLuGABIQS7jZUsVWId0Dq
cCvh1DvW9F8X/dk2xAYH3AjTa96UC03e/vgkkQrvrEvH6V8Fis0tBnb76MzsTzKkWMxEIC4A3+h4
6916GRhaS1xDqBUyM5+WFSm+y/uFKRFU3xBBAckqxU1l3hATS0eO5jhz9AhjqB0ivjB7H/6VMa9h
clhQJVYznNbfpwuQIfhifCCfQ5pOJjbSseUjToQ6UHb2RIv5lVMnVtoOzvWVo8DLcvoOCniRysm7
Sk71nN2fSIkav3IY7H/q4U1pgK/7RwD3XI7hP+GrhHP5pzh8YiR8IMzNGFTTsWe1+TgJD+bZVR8H
YIKqyvVVvIF1I3N7HafIXKCxIFUf+s6JDUy6KsIP94F5qres67kqLoaKx9yODHPKREELfYnkQaLC
6DDJN9FLUtpLcotTa7Rppj5lpWGaQKzVOV8J+TcRnrR5trZ1nU4Bdq2sXXJT7nNQuv/bkBYH7zvr
F5mHJn2tAhHdBVTtyDsA5MjgGGtwICoQJzHaO1IKssnLVHA5+pwQWgutFnfDRcMeonzL6u7vLf04
rmH0M54HZMrjnsEb5qNH+WscGDbxMj0g+Y7tB3VtKIhobNNiKAfIX7b4ZI3EIyOKbOt9d4BMHDCp
WHU+JNHGPTKwoTsB6gHdccLjEHoUlL/4ZkVdWeRzFBrn91suqlrIVDga6vG9MG83UHpA/uytYeta
g91upNBslsg1ko13AXj1mXZ1RYCmqVgGNe+U+lzzpaermBZ6xxZgUXbb9aCm9mFqrEs/gj583ncU
sRYxsIy7s7wmwzynwVQK5bWTEeWTuglXN9TDVS1RXbJxd+K3+X8LOCkfWhWWXJuoZMK2DYYAAK7+
1oSsRqSoQPgQ5YscqAhiZbF+Fm5ReflocYUOpNH5uydMLlHPVZpnVEw1LbkQ0j8gqctC0DcsSfRP
mc+rQJNgxuiODoa/VkexOOJb44ft6gL9MsSp/MmmjajaZ27vFUCYaYhhZwPiIG3cLu3a0K5q0XO7
MTl9ZajUqOdrXBxsUwc77nXZzUe+FUxSi6EZiwou2X5OY4dSsD0ZKDi0oVdLlDdY9vz6b4rFNwH9
jM0g3NQisT70SPGAMJKRHdAm82/hUul6CJGMxQ4RNvQBlofoJi02oRY5mSDD0hGvfPDK2+/2SirC
cAbUfmI4RqEzWXlgoEIg4U+JQ1xxyBT/q5RvLnAGRHMdSbdDMf5VrHrHKF5CHrDNxRHJhcXuWsjb
X7loysx/KaloYtcmrJczHw1oT53KmGqsm+oe26fAGri1mGWKfUL1j1fMIjZMjTnolWolfKIRefvA
DWjrjD+zMrldwCmb+SH5oaeD+itWxARzoPm7Y4nZr2iN9WVPe7cAsYejOWkEAJa8/iD+NbQW8bqd
0Wkb/6qmdBLkr9Qkh4WpIHKTDRw5IFl4Ng4K62D3Ie21NihvjPryClHp9d+TChY4PfupXemuprkU
8xspmoXPzHJLiuPck8uPkzrWxP/T5ISjBEKw1UFyrnWE9u6r755z852JRqeAz81Ft94dwzUFBhrH
AQoCLfYIkI6e904DMOSorsJm6O7f3JFxZP8WLbTkQynnvSQNHQnersUEmPSmiuM8nxqJw9saz19r
Zrv9iECOOz+pQz6nMiMHVmxf12Qr4T35P/eosLsZeaDavLEZbSW6YIl3P4pnhLypF/EyF6p7rV11
tpPa6sgutLiaRvtb+uIIh3T0pASKr7MNfZL+z4R9XuuHmdlX/xPsr75AIB8yYjB4KsbKO201GyGh
TtF4jU6PV5j2uWYvRBWNNEdwE7H4Y/RW+xzfIDT8RHH3AC4liYU4dK8/gg1xvGobgVmmUZNNEMXV
NGaRPccziBDMbohmDRknU+dNHRjKhuimeUCAFPDJuKcgg2o61hk8zgvKX+zqs/ZjQ0Bk1WIdpmZp
FC02JAL4gi2nkG9RCdEJI8e4hQya+7YWc3QhFtQhk8/SOG7AzACjVNEuPn8DUUu6vEFwhv5GbVbI
shkthrHUYeC8cyL+1xh+zwKcuipk/gpmYZlv6hn7m+5UhwMP/1w7ItjT5T4Wcp3bYSAA+IiV4vOr
Z46y4qDBzctIeaUSx5b+/eJQ0kwMf+s5P5UIX0QT+iv0flM18Gtybz4jK4YRRgm5Cq9p8xpSvA3O
vdWiCtORmLAu9OFkFAMagBa+HleMKLF/1FckeGUsm0dS+r2O1JQVC0Q9bK3p0iyWYO6AuZimTw2T
ZxQ3xSXNi09RYtNGXyrQC7AntH7bERHAIv37x8Sq2H7AAHBtNNSENghsyKRB8uKN6+Zs84bmJfJN
xpbNrRKAOYSBbU4P+vBJM/GLou/5hz9UwvhHCh2/uSqwPRzhLAcVy8oxEYbMvo4E/NfNq+t85+g4
lCMj/zauDCoQOAftvGqM4v60eF3aaODCPJzQE8WFBtZzMIAhW4tZrki/sQn2zOxjWOsm6Ib8RmtX
aO3XIaOuwxnLuphs/Bg60Hj9u0WjYaeXifOddRjznSze2FJ2w4hHBMd+UeEW8gSvW2diSnH0p74f
yaLWSbPHVC3HUo2161tGgLWdodvZCUwhrZYSA+E2To0jOoguI2gRgwjpfx4MWBD3TVgNRtmby8A5
fGdG4rAcIKiigIyTr597h/EyOUUxWeMdPmFlfcPK5U+f5lNf11nWZBzvVgW7K4NHcA8ECxonxlxi
L7eF2i7XOaepycHvfEKbcMyn3OQkEhf57Boum+b/Odzf02c7PUScYjKYDk6o2enHZ3dXlnTZoRWH
D7ex26OuSf/VipE/qdXGXTt9nubkw3Y+tEUX9MtxZy2kLeEeUroUN0NoCepdeimPGa+nTBAu2kaE
1hn+XWtjh+rNUdY+y2e18rZ4xEkoAYL8e73/6Noj/mG4CSPOKKPAIgW+9SdY6vNBVjR66+w1zHGz
6uzGcUZJOwmSJwiWMh8Skzg52x9I4v/bVeHxph+U9ZNQAuh6CTqCpkw0LoCaEQQmbDN5494beQj+
512ZV9oYdmLcwfOLTU0Xh3PtgLNlcK5STEBbNXAU67p4YvevJg62SSZnv+hjhuX7xhJwX9gaN8eA
KoaTBR0x0zYoqLVT14BLaJaYbEBucPFFri4t/Ie02mw2Wz1UhgzwaLdRRGAJLr/Hh9ShC/T3CM4m
uzicw6o6z0iZ/nFefmA6uOOw5FBxBszdIf1uxAyg2odkRwF7HNW98O18Yy18JCp7Fp8sLwCpcO+0
2ocro8btJhK4YiW5rgDhA51AWAYysJ5z7AkImqb6GgORRAN65Jfaft6EdhtM/SdZ4bbmYFXmPjiy
5H/OeF0qmS0obZbqVe6y3QK15Y58hv5oNxRb+K/QERLeqz0swsXwrGoot0xiZIH8SoaO7Dz5lbXT
r0nqsbx7LdvaUO0gEIRwWguw+AVLasSGCqJQmRtF9IHXGfEiUY0ZBG2lKEdOPz8j+MJaSWzhMNNP
1N5G4hkgThD8otB5SCGK0zB39fdaA3Q2dU8inarUDKB53dYg/cslt8/EHVROhM+3A+ybf0hx8Cb0
jvqNo7LioInmpj88Q4psW1lkYd7AFy4LWIdiMwaZvWxni/4vt/zhfnqtJwkh9PhO3rn0zeeSVahg
ai5KMzHjCXkesfKzE35S6hsIjrRjl9DnA/UbOjGkcSxAL0JwbwLB1GZb29XWUOEf9fFUMuNo6tmQ
tTLl/OWC17R7n06lAplQqEHJS+yEyQYIGEMVKMGvrYHcPyycMhn3F3+8cqsWswxNUsGsHNGYr1MJ
UsQ0ccirDKJY9hQnn0KVZ5JCmcHGD1t5cJUCH6TW+vmaLu+BrM+DcFHYoetKjMVNN6mn8mkBAPzN
9TLnKod5YkxhIEt1hjmuwKcdPEZal7IHEBPAq42UM7E+T7Jrzx2mBOCG8K+1levNjnRCr+ngSf4H
reW/LWQpA6qXO9Use4al8N2UY3mkLPeRHWAQ9h9Ue61iuLb4wlngmqCBllrcNnyw22LsCQeLPuno
o9yjyl0w3DibMxpWcnQWKNiWLfk4K2HpzonDPfQP0rI++fCgwMWHkdkS/iFY9sQOZAZ9Ks0NocH8
FxJ+q7T5uXA3jnXETP4oNEmOo9Arpd2Ixg2cyGEE2yPxN5mhawNvTGnnbnDGvF4u++821Y08iMO3
2jeupgIeY71T8PEkkWLwdNrahRLZA0ggXnVBRxnCFm/L4c2xKlUu/2TeFjXr6YpCWRhHJ61Rozjt
ShaPwp76WoHpmPtZSIG2f4RzXQv3HGGyyWP4D8/DU/OhD0qEKIOUcOH04742s+5Yw9aVtRNLGEkM
BAHxmA3uH0u8ai0Z9Ox5SqRfpjeFMlqCAhX3j2i/5dga0cjFyKY1poWJ0c+c7kCF7BlpG7RPYJbf
NQDxLs9hmD/N55UzcMwFVhaqBkFdUL9q5VV6W3DseltnhkCGox6u+QW7zprY2aOLM8BW9IbF2WGn
C27McpfeYK8u1jcuKMZsmPu3HRkns5X2l1ixE2emUXyPTHYnk1TI/GVg4nPeJN+Ndl2H1MzcOotN
BwSlYZaypzEmbYxKQ/MBOV2WeuiP/dyzK5p8WtzdF3qNbp5jYtr80Zq8s+vWRgWnk/FzaDp8AzR3
AL0+NQgFP55vIF15OBq1VLkX7KT36nlyIGDvIvfUsEH/HiiX02MTZKnvJ3Owx/4a4p0O8UtkmNoS
s1SWs+9h67e5LkBcsloVuELuOrHxuDKwtn+Ne0bZEEETbhGGrfsC7c1t2I6rcu6PfNtoX3Jw/DQq
pWBqu3FmSVKO5KJJ18DYpnSVbX2gG8TzeK8LsjGM85LPoPlXir5+I6hDpAoPcIxcYO/nW6qNl9G9
q2RWVMt8c9d9tPyY4MoCJb3Of1oGwEh0twyviqgpxBdDVPW/xDIz10j09jKgoASMpIKdP8uHWUet
bJQvKIH/ux//hNYpMJFIGbdBVsXRQxIvI50EAkJ/ekIRBnZI4rDrwWWFLOhW7NxgAq1S8mf6msLO
ah6M67bHuwDfx5waaTC9Guoj19Ba2vqThjYv9xcart+z7JZoP+BzSCn1n6wu6F1D9Mu3CcpOPujG
M6Cxkj1mfSfsVZUO+gqoUKRi7Zjm8CpTzp9ARGLRalqs8dUUL6XHq3CP+Jxoy0Ip2kUMGapD5zug
m5m73Kkp3vM6zTX6F0QudWpDUgGD5Bg+PfHpxjVxTz5YqZbKNBNeiAUKwNUreTdr8dRKksEPCojq
uc8aNahq9BwUjRI9GcPlmLXZwUON6hF3hYwd4atGNU99ZkEcElrcbxs0kl8mwzTZwe5zPi0y/k7y
PHAHecfS+K8PcMHAIx7JTn+ICnWBvZLR4F2ulz6PGRIrb/ATinpZk+ykMbD/F63M1X5bw6BQSo0S
9T2h/WRMyOCNaGFWDry/JTQdkFCONj5b72+sntEK+afalls0XzyB4VnK/ezlxmweSqNbPGxZhslh
XT7RjU4CpEVnkPgdBSy7z2RfgS/eGGt+9a4XTrX2hoW1xk2ybTaKP5udWCWNoB8bLAznq3f1lqyf
rFbbjYS3xeKRFqBjRR3O4KGEcERJKeQ5DAXDVGwOuevWlofCahVDPym6XKTXlfaSvMrx1Rn2t+h+
0GOEbpCui3quLApsCS5x+y3h1GaVXTkcmmOPHvzhwL630z29fBQzQUSLknc8OwChejxxlPjSXV/3
GiZq3xfzkj4FaWjVeEwc8G07vM+T7Iu7Zq/ZKApkBvfd/BY8KpFkjtcBgzNoYiy2H04XeNzdF4Aw
HWMD4/d6LZQHVuXGr5AFPyxAFbXngKFbUjk1bol5s0cLyWVDOw1ChgqHiqSMtEVPaFM3R72lsGM/
vYfzf8//J8rReJQ3n9r0K6lFka7rreYsL6dZnX0O0xerxeqhKMKz8pQSKfVxIK4wbl03NxnWMBi0
dqSfpZE57VNuem2/6lZnps2OUnO3vzSMAXvyQvnNo4hd79ZuHNtV8l4rOY8jE6W3F2MkC2DClZEz
xkYbhZ0k8UnIddfYlHnA37ooVqzQxCSJ49ZXXZ/whr9dvD5EiTRHMLLCwPZ0Y4MHvsbfzZUXVCAC
D0ecvUeZIcOwU6h6Pd8Iqfbf94jClwa2ksHx/Z9rmkgSsu8vrxfOGJQ3zz/GsR8BNad3/70d7G68
PGUPET59nXb41WCQRBOGSRQGkGOtGf6pAu+67E7c0CGXqP2Rpky1Y35E5lBQR5mVy2ld+JX9CwEv
7CSHtzBFwXmr43IyUpVadleUeiGLq19u1M0dCXkDpeKO97pIzlDfbvs/nC8tc0fDzPF90c46u83a
2+W9LOXBothJz/70fy6t/S6tysjDZ9FRFOQRxMDbJ6Q+4e6RWnidatc/MNRU0z2F0f/QYFbO4sYL
FQezZhNN2BG75xxAfupvq2lS+8IJ6SDGjkQG698Dw8vMS4POTYJ/4HtvfwNpauHWpfckOvdM2Gjp
qIkA8JsCaBaMllIOLaJzfssi+8+Mf9q5lxde0p8/MbxD/jXyoLiJbLpTJ2QllY1oWfejnJfXY0Ye
iEJNfjjseqICEsv2ZhRa/psBODz8YRExAIwGtKFA8w3FlmPkvrkFuDrZDo36GlB9hbqQyTwf7uIP
Wt60kwiHrObIs0NdfR5IhGrQPyJGjlf7ZJ+AwknHGV7Mmuq2FsdriPzcCIlL90JJgOlLs/Rb+1LP
lshDUyqBOkkla5uU4IYJjmNcpu5zqzt8DpygNeI7YD////A78IQxGur8SVt5iJJSYUZollycWZ8H
qNfHzG3oBeZfoCWWQ9YS7REaxAWsNzxdeQtEyQfBOV41ORLDCZSQaQX3Yx9Ux3q6C7bBpaf/xN4m
JB0pXIm2u8wsnn6VEFruQGPX7SUUUr15o+Tq+1A8qAP+VBp2Ae/YY5MQCp4Njjl2Qzn1cGQFNs1s
sdNXEqTofWrsyXW3y8cStgi3NRXX3Ol4feYCZA9vpnxEVcLOqpEPotZ41bFEPexRwoJ6GZHtQX90
bNp55pCfJnN9gm4M+qnV7y8vTgx897eKABrNy/7KMDm9YgNSttraRaYeUjyIxDpj2WyovNt4XGY3
iCLmskzZWu461N/WpjQkK8IRAHzKvpgNCey7E7uS3rHRJkv0Nt/UcJG4dad4AfNj+xWYKgchPpV7
8ZqEGxoqHqapGBdwu/tRdZgXVWEimm2SWhPGk926Jbzmtr7Gz01iWS2iLubNjWjTbOcEITAT/l6P
6BxkPCI7HfXLpgOGkPTekseNIdqb9mCQzqce6U+2ZKowhaNO8UaEGwJNcomBqMIvA5ANmgFy0hx5
BI+5OVbIySmfAKn2XB0bj9MdfDjmrzvuq1wvxnqabCbDXzlBkLcd4gv1Oj7Q4OXW99Mt6w6ATcC5
E7ui/qCeBYlY62cl1yxYKuLIRzC9AEroYB35LAtYMlybeiQYMg6rp6i7AZnOu5nn8HItWy5q6B0n
b5pBF0fOIwcYiA92bEaVqcJrm9KBs4dVlwFmTNwbhrQGVEphcPwgI3NfA3h+Hgogy8xtayHEqkR3
qnsKa/ex8MYJ0CCpVczA3DiTRCi0siML96Ph+PlukF4z9xdivERyCyaRT4FykSmNTMt9sWkA2u0/
/K92Cl4AJ/Na6IgMeTeLkY0XolphpgfcYRH/mXBgrPkc+rmq5hWYl1Sg/CtJauGnjGHerxkPrAZf
8kVeNjvuiASrr3/LJN/ilFg0XrTg58MjcV2phqDaOsbpuybC9xrTLnpmsjIaQzPTcqRjdPUhwyfY
1uWuM8tBIHvIx+H2P6RD/vDzrEGo1KQJOrRlevfz2jbKbn16vSJ8kWOX5UKcGdyV1ryUqbuHEX8g
UxdqZMBpQHcf9CGfgtG2UkC+3hYG3EGlnkymbZI8gxsfeWgDVP2Y9XqbwBOQgthHIyyin0eqKMQq
7bdwy1lLQEho3M6LyccO3oZKQxjJEovcwNRH7SNOT2PCaGGXBG0/9rzcvEtElJIlSGm9XNIciv6L
uNNt03Cw0EUwZUbh2yRcsPIychGedWlhUW9fPBed1/Q02uRFfKKU/bMmI5xnGE9eoAFur2aYow9s
CYHNtY1GS7h0Cou8xIg7hoUmCqo/tbmM3RjnXh987d4loXsuAnQMpx91ZgyV/nvBpsJsUceiE500
94ki9FTWyoPX1i9O2a1J2K/n16pB1TQZgXB/McSCkSKQhbsD9fZyIVJAJj6X5raRcREtreT1zd4j
TrydanSWcRbi7tAeljM3iRrhbIugAh9/lG/2QdV/oUwIudbGkI6ZAV4A+nNMZ60+z8BCWjLj8/P2
G9UvzlCjIXpBGtDwfJZ7XLcynqWU1MKU7vJk3ThaUcxiYIaqpqXvbKnxdtsvVbM6qEC0R+6b1YT+
4x6i2rrJnvIeSLs1xRXEF16el71iAxx1Xr4c00vfapLaWdVQ1iosYX4iNqKjGUWGKgCBms8kTQmz
ASb/J0puVsLZrzdjibbn5chCSAGryxJz25hvlwgXJwpwMGmG/hKJq68FkE+xwCY+WhfiCyL0dl2u
uA/OcyI0hF6MPa3dv+7kru5QGBk/AMSOGyEqlIZNxjLm0kDA2VLZ4kyN7I9jscnB7F/Re4aECHMA
VvkJ0qpZ57MkUA4BAYNmBzIRUK55bVsRaiBky3YdXvTUBGHtTq1TEhgfYyCLaT5q4OJUugR8cWRO
ya/J+2U678g12sWeO6K1U9VU0v8cXjb0J3DvBlCDOYP/ZPgbwOaDOtqqHmAPvGxtS5DYgyoeD4hr
u2RkNwGZ6R6Uwt2lFOfb6E/ZHOS/E/+l6na2gugv3dmn8pYISSKudiamls5gHQqWCo7lmSE4TcGz
TbDGK5I2hIq52r5EY+FADY2qlFj4b+84XQvKpTahcUaLOohgNCXy4RIXpc6MJJHJO7T40GlUhWYp
fp/1Y5G+45xa81s0ZOePPJ7WXoKoUbwp+ZcW2Az2BhZX6ROjI6k31CEEGlUrZvV1dcmQWnOUi82t
fPuFz2hdwIfENYUkQmlX4eKND3CHRgKTLH2bJYpt/UJE2f+SjxOvax3YA1gABvzp1HBF36zrUHVd
hlmwZ0QXVjEYoSnrzaxnNDFW6sAO7WftSNk0I8JJhD8xBl1STgNt8Tk/All91uz2ZIFrY9S8WaeC
1hhvVtcpsqIVVKErgR6fxS5OAAz4mExj/BpD2dG/986ZvYyoWmz/QXYcpHzHthIUrP5a/rtm58CV
3eVyNedo6dhIehoTdgE2HO/NyhJSuCyGk/n1dfExAdY2zWE5Fc3ern0zxwgDrnFUNyo++clCPF38
sZfp22yBQvZlh+oazGT1BtuBQEsjotQME2PdR8StLUo3Ou9WAI1/sorBHngICwKaEUQ0ATKQQYnR
8sxb+Z5/bGSibc4d+EF14l8KZzTj98G2EH3i1gkb8OvXVrC3nTP/dMPfsj5jGGNksp3RtFSYTtUL
SpY3yZp8Sl2vP+PDqZ4PfAnITXwbr1rdXl3lblQZCW2Qntsxa4qN+bghzf91E7r4EsIqkgpCj6fL
Q2/k3Jqw6hwg7/DlZy+cKaoF8lHh5a4FmEVXLFHLDjh5xktWnkGe7I65yTn+P2N0tYp0L6/q9yyI
/UwAUyGa7B0ZFo4ExJWXvyWINAl+ksZNWfMC0bDAIh4QdfhaTiR9wQbfVwElB3MMBM3KTBmbFjJp
Lw4MWplOM8Y+aJK81uLVP+NsEJrIF+iBMClYSuoF+jOXXPM74xRiULLrlSl3nGr8zQJJh+QZHvfv
lKnoP1rWxyMDSEdP3VrssNdR+rhhyBHNU+m6DAwfYWhh7larBgUr/qZObi4f5CiYf0BbUOYPgn24
aMY9y78cVDnYXPLg0WIGULEWUcPN1beiaTMt29XnY9D4Tiu6plgVWSckxScb80G9hLg/vMI969d2
PCf6frpnLGiNTznZ8XNinvGX7i4WOtL02FMLWohw51U8tP9ztdzehlv2AWY8F6nj10h4dSw63aIh
QaV8L+VQ35Gm2CJrnM5lkRJfsGyIZqUxwWbH8/GVmT7RZNq8SyE74bybE3xv747nubmgxOp860v8
JkvEXhqBFa/IhpQTUATE3UV1iE0W89JgNxnhtSJpQc5AA8vYnWkd3oZ98f8Af8DsgLHR+RnZzqp8
vxmu8rovJH+6NQPxdN9OCeD1ot9uFB5z6LivSHamuXIQFCPBIBUucNqF5v4c1bnFcIDMmaLKmYX6
k3FYJ/CRDIbJ9b24wsxbjtjrlnx+qF5emyM7ZePHxIDcrtwT+5KpclOQN9KiDhQAUFNZBtemey7M
VkR6GxFD4qr7m4UPjiQ0RLbUKfTQ9fi8KAfqTxaHyXn8Os7Y0hOnVodiC5tKW/34ccpFl1ysEFxZ
+jLW549Or+mNg+a+RTk47y5lCh9PyIZ/FyqXFTx5dMW2iPXuMCTW6fTkpJdH8uPCXZgGcyEXavQY
savHOi4VrFS8wyVIhbwvEVj+ovyMYkFQJQsrmA0oFxPyTK1ArPUcwrrRrBZ7CrQ7kKLABRxXelbd
KrZ5iTzfD002XK/XDHv+NeUez1GWrqwUnyHxtPR/JGpweu8dcOuqrhX87zQe4no3Cgxu6o5W+HJ/
1zgeRSdMNQOXvigTzUc3VCZQlf0XR6vsWQC3oMKZM6FQdCf1gvhhi3+eP0fHIHDjwQwxHFCxQSNq
elux6+Cm4elkOm81xvC0YPWJCZfboyq58/OIPbkzmzlCWxBqI2P+M+pObqu1qrBYbcEmb63lqUQp
ilIyGLIuPC30F+yP/vqkCS79bkHb8z9fjMnFLjjHW+losrzrhggP9v/3u6BKjdHPrzUT5I54R+7j
AkbGoX+ikd4Q92MsUz2gz69dzx1/BtRAcRqvG4+S3F8oNzF4879hNVPKf04JMOsFFmGJbG7zQhkb
04W7fRmWkNVswy8jlAAXcg71gu5GLgzn4bx77x7fj7LzXOPzFEOUXOtTIAqVnMNwAHSOjWYoRdom
IbrAXZYVFSnm13rh4HOaSVAxy4m4yFvTt4zAZurypw2Vc9TGqrqCKzWhjS+RAhs8hM2oY9TxJXMM
vPY72POXE1W2uwfMUR5PWHwnyCOmF1lor2jHP7Z3FayYLDGBRJp8x1D4y+s875HOC/cr3lm/uL3V
oDI3U+vt5JaG/FwsXWXz8F0XDdpXzipB5w/86eRTS3RKBDPxMfivb13wweugPQAQNCZWdjnxxYr4
wYefpVQKYKPjTM2dl5CDcMuVZ3VULG8UE8kW+XO2DW/ARqB4znoH5NFPgza7GCO7p/pwrpOX9jn3
yH7mXM8wL8KsL13cD5mla0KFHt//OAFhiLOoRSGI9kF1C1que3HJucGLfneH/Rm+9nVAnCI+uy5R
6r4lWzwnj/++kqLhmBN4lM6KaKwrlt7fUq7uDhoEdJZVFqwD0Y5EuV5KgFfCB311yR+L2TfHee/c
zNs+TM/fL5tf40DoLWR+vkbJV47VI/bDoVxz+D5RET6PRx5BRNEg2IKVG1z6JauzKInlBQaoBgkD
g3fhqiCrpWR3sTiMUH3UMh81CD3JyvezWz73ERrv6IzilQSqb5TwV7I0/0tlhZ8byXVyPfFdOJnn
hsYignwU6SrWQS4l+fC40KC9Fs5aOeUifc+CYxmkX4vj2+GCiGrZM7j34PrrXFGEjhbLDmkQaZVJ
gVnJt+7V3eoBlx5Byl6iWKTZOwQqK3VjsJznA2btZh96dAfDt43oAmLOL8ZCMECCwCGXylBS4Os5
QYtFgslDaomD0pgdzvKKQ9K5sS5pR3GuSuvad+KBS9yMMeRc9iil3kSbWJ+gQkeUKcgxIpVgUWSJ
5X7ELt+/D2eFmoLxPScbAfIgXxHFBu6PuTAohSP96+37Iz0RUSXwb/ZQ8+V2wtjm8y8JxyZVqYyo
NETioQe2NLjo88hyT1L8e1ZFh9oQpyeFlvCY+zCYRMGZE1r0dTgAL5HndO0LrWrQ/6g4laU52YQr
FGFT/kJnu7XhSryAyP1tle6R5HC1tOsKZwIhVcCipUInCYk20qheVjHZrEurhCkkioI45/Uz4Bo+
DgtpFeHYZ+rL+9PM5Uf0n3zum2Hw0HYLculovsGd3UFtx1g0cnW0+F/UjkuJUiggvPCCG7SS/awt
4Uq8AchHIYlJHjkVZTwjuyH1uWpp9AREPD+SZTXjDIydbIPwH7zvUP9mBVal0oh17w1/3vphyBhc
dIUFEt1bvAG2KW5eC0mjz0DG9Ocq41d4k5rlEOHje4rzRB+vSHL0Jja2UieaT7iCg8uuN7T7569D
4MRHuyM07sDrNlXsfR+AOWF8iotcOVtpwXWN2hvvKudODlWc1f5CsMWuDj7BwJKmfVKNnLNPgbF1
c/iXueAlb6Em26KntDVzJy/vrCnRYc+nemZE8um3gl1PmKWjqpGlnblBlBpL8HSESAFjZ9QMlM6O
eRz382Yt831JcxaHPUxi1YP1fQ/ug1p67vGT4EJWJTBrIsAf2NKScshsbNzoxYUJ8f8wIIvziqrf
unAQIlYRPA+f9QRtVSxD4hytik7rdKA6y7eErjM5SHVkbzsryEgu5TE7nuF9LisbHVSrR+8QlUPH
9lpnNutfzvKrQQjyMcwepPTNXL89MyU0sonhpZC+HtBadnai6GYmecXh0V+T/Zcf8VCw7K48R161
nIMD7nRYXfMxZLFna6gtFel6gFTLda+uiKA3ci95FdPij31NhMK5/qsBJhqTNOdJnnMCJp7H6Ofk
NUHj6cNZZtftMkxTPbm4LtI20B+4nxQwLnhYMPbT6955bVmFVmaZSm3hVNO3RXneRLVl6tQdRJKk
fuieOpJoKBFMiHNjU+1kyVtSSmU/KcDCzJJFfdnDz/mdFwM05aIbIRumgywqOAvXeoIwXSp3fhxM
MzcYIQ/jwtkg8p1DBuxR10dfh8WZOtwpg+/Ati+nSJsRQa+rti15gV8RgvaDzlZEbaQJ9o5pOdPZ
66KdeHGXrNrXRBsvHOtuea5PW0fZ0vXEspDdKlpwcAammIzqOxJ6vXZsz+2osSpDr0/d8N863Ztf
03VnIptGE+vzeWAuJbTTguePdmXbV1lIX8I24RUQTNHauTvUzenIjDYqmTME3+7IbeYRE62qNTtJ
/4tVur9vCQGgtw/42y8CxkC9APTQc2t8/ccbSXxIelRHAjibDCNGGKNWsLiGz49cDku1jNARa8Rw
wly2v9Ce6dB4owhkWbyroZZqrJnhwJdDsakeP5f3mXWClbfaTXgHwJL/7NiF6/PofE/v/OMyRjRS
e7jC0nAYlhuoT0BnNaHhGvz53DM0y7h/UKZsGaihnNkmHtjSUlKc4Rt33Vhm7Qbr/ldIVt4U5Xhx
EubJPcp4QxJkThogk84s8bP0TJr76vQ1xlZMVa8xu5AVVJewXvHEnIOgL4qyk1J02QN8fI9DFu3d
mlsV9L1h/vlDoJ7G1snCDmLFs12mRpg652lfbmUMjL8sZzOUpek60WxC5FN9uQoZlKVj2bD9hZUQ
PTVvu0BMu0ixIQlVrvWrLrJ6PC+HREMZGHwukV+oSgCtTSALSno5LYRQzH8XeYeWtZTU0uSj8svw
VP5pLKvQ62+HArq3JCikWc+iWlPu7pVhTfwWJTxiQJpe8RVk0LutP7pD1HfUIgw+xzkl1reYN2Cw
gY3uBUyXn0h+p8BdzwIc1ReXhwSZifmQxmtkTHALmL72SJLjKrHnqazAtN2hMYvdwG27y2RuNlvH
wURNtSEs7SREQSFaFkWAO4+qTSGa2EUBHaWvq+FCebGYocuIY0PyP7MF1TnbZOzYC7NFj3D6LIDB
3MJL2/45O92qo2dmlLwgERZCK+cw4z4oNAyCytMhRwHbxuRjC9vfpTrKpjXjYL60+LJuK+h9ulE1
1IiuF2YIpBVWgsB2bA0PFRbZmc8H8EJkD6e+ltu1Rc2ZAViYd03+7dj5cNFr1AwUiix4fI9aCRt2
v2BJQd8x6ODFxOfQvUfsnrtC9Vkg0v/T0dbZkI95oeITi/TgCkEI0poYy7+CekZWRGfSu6a3Fmy4
eYguEZzeli869IDySiv07clxqmI40jcrxKgfRR6O2ukgmZ9VlVoQwh223UzruhfccCittFxROVZl
Hw8NEq0mukzorO9EbSNRiMqz1EUq+M+D/hmWjYgpYcTHdjcTbad2zhUn1lfRNpWOXspuYrEvPD/q
cT49A9hIYVzkd0cKM040Emix5IDLMjW3SNrII3zA8xe7qNJKdO9TQC3Ry0g2e5OMUqDDjSsMk/bd
98urDJOK5tdUzqFwCQYl/2+xbCSrCCfu2CFPtbCXbdRQtc1ImAfDtb0R9aVAcr2P3JjM3EvwF4FJ
VOZyyp5my3hhcySDHmioFXakpzuWMkUwmsOmcB5rMxfmwuYOM/2uEPYcdJ94Bt33ZCa0EiZeJJ19
6HmXtUdINtcg2pth50QPmxPBQM87rC1x9zJ4TRbFTR7VsC/qQrQeZH0v9rWDlMxiDy64/yGm4ZKu
FVcBDBMhX0Vn6r0cO+9UaKkHjjRYX+gQl3Mj5DcaSDckZsaJ1ZfLmdwaxf5iK/S+/e6gik/egdF4
OdKBydeZ3olSGHprlMqF35X1jAitUj+ozoWHVgkXD9ce9qfCb0je9utVTM6igbHJ0j6L+lAbAcNe
+UWVopVAl1EqW4Wim0bNKMS7tjHGQVYXXjBpEnfdHcu2znOtO6iZRgDE2qkhHbYFDsRb42mkf9MD
7WcrOGo7QlHDGwiHcyPO24Zj8P0DXMApnzXo0UrjLzX9HVBR38BIrfM27UGDaTw2xMHy2qIKPNsu
M8w8D8aabPzFYmUaJyMQ45osCB60L8o9ukHCBwa2ndJhY+QJkCb9eG/hQY2EOiy/nFLXJxgzG03+
VLJHnC3sYr3kzH/A1ez5gNsQgi4HLZRNnGIUo5IbQil90O7w7xTFPYhNpVyIaw9PvasAlMrZsRbX
dfWWSj7cXm1F4O49G00cy8A4MxZty/eixqwM9rBRkh2uiq6vZQVH+UYOEjktFv87I5rCEz3jWtCn
bjOVuT4oVFdOm40tejN93Pik9Vw19qYIhXTOKqltYW9tJG9z/9sZHhnynUt9mVlJDd/2C8BF627U
r3XheJwoZT0Q2dl4DiyPJ14ecmUiDmjHZlK8tFmRzDeYeXIyNXzo9A05NPn6VPiBnTJSYiF9APdN
TIlANhBz5lYqNFRTm3b0GLcqGSibfQ3Lxz6SSH0gM66lKJzmTdo8xgZfsk9oKpw+IoVhIiCVJgHn
EDN1VP5pYsd6zHAAP7PHTHAyES9Shlu6jeVHpL7VtQu54/R9+NRl5vsojpjoKGW8GlYcpJ4YefiE
+uspFCSNaii8384DrVflRQUurTEPBjqdYKBbwd56gmJfDpp3czgBuPiSuo5TR6l1Js1V5zew+tlY
ghb0b6ja1qInNGBKNOp4y2eN1QY7dAJTDatys/r5RpPA6OFNTMWeVDzfftraTKaUHi4GgilzUZUW
7p5ddUgTR2iEZCcEFFJiMMmUoo/AFEDtztdkUrt0IbULosdLCxSb4oiHoTegLSN2BhZ554dsIzJA
EigQB/CeDNsuPaRdYjPD9x3vHTi9UrU5NLQBsdBwoqSYPvYoeWZnX+lHI8lDec+/Pu93pljiP8B1
kZLpb4WyP3Yxrpb/S/oqEgbNa8IfUsYHgGNuYQsBj/atDnIh6U67/lxojSnr6w9Y6J/wY++Cuuhg
f75eyKG6QSR7fp2IzZ0Mr/bIvq4Ieb+QL0klMZx4x9bUV6ian5ThFMtDJjISyaYUdJzO/84kz/Zd
yzZ1NdGUckhZlHmL7q/CWlINRk9QjctPOUu1xuuA/tcZl0blf8TMNgaIadOOTjY72RxkrBfDw9tR
nrr/mD+Qvil04z8AfUqgjfKG0wPBzbTsBOmysV6Qik9Ydqms3cKZiYMpHjI4dw5aKX8IEDuuGpku
HbmHVLKYrCdCaRBbBEe7Bii6U6fY2Vd7c5glCoUBurCCMoBp+s88Qa7AHJ2EtM7nkBlXo8CbRmpp
UM1ayC9GAb+9pJbAk5RgyRM1eQpvIo37wSsXpdPvN/oP5ZuL1tJqWNIeZuKnyLHN3NFyYqDQxFZL
IGEViRTYajNEEeySThcm06IfkF3ZWAlcT7BB0mJyXE09EvJnkRyu2/UbwKpL/SBJmO8z6LvM5VkJ
T0i4Gxo3HS51nfx0hkdV44FZQCm0aS4qLoCjXRkYsuEpTw29fXRE6rvJJKwvSI6QBSdsnWvxRok7
qHdECc26X+f0Qyf5yHR8CNyCZGWJJtrNQE594E1YBpsUgm/vG4ld52f5XOSxcnsl9EItj1O9o5vi
7uiboofLDiE2byNWrkqIYztzOlCvuSEtcfVMguVHFpzSP5piJqRGsuKmHjynxSWj8fyQe+sIHp9I
DnENU2BowHo2Qf35EbeuIQ0fdlv1DrCZpY51i1/mIOjytndeNU042fev65T43quTeOSwrHm8RrOZ
Vbhb1hJtTt7B1GnXBZd47+AikNNPEQS8hmwO7Pd5j+OBEgfUIn21xeN+eQoROeeEry+tc+BGfsmV
e26WMg25HXD3ZHDZY+EhWmODEwcXiW0KjBFvPIKCnL1RIg+tYf85WOpaKn9S0+mutB4hr+x6V+jQ
HkchdFrAFkN07JSoYojWNEuEGZ8iEHvIv6bv3miMjuBnGBArjpM4uKknuaDlAheouBnK5ex170VV
1wmVVRlQxecacs1zTk4WYdC+cVOb3E+/P/REakCnLgqi6aUajeurszlg2cDwzGae9CpDhPU4Mroc
+uBCi9/WV7JhBd4idkPddGnCrcrxbdwdmX3LinihZXqFvzeZ459RIKbjVaS1LyDynRyMCFoiJjWB
TlzN9iZR0juwKD/4TYCbkLhJCVKQBYHyihFSlKZD/l6a7Vwo5SQ3bf1bRkv1as9TZWLSdnrBH8R0
BNs1bUbpRJRD71Q/8HB5qBh3A+2YJKFFBqu+e8djMpN6XxFwC0PKAajMhSKg/wRGu3Lzo3lq75lF
6tdwM+kP4RT5AxYLLMc/CY90GHLgnyTAeoe7Jfmf07o8Z3kWlfV0Mq2JmAYh9dpUS34RdYNJd3hc
JbRApb7MPYDZpqiLHbXIYI1/Ai/skMQ5mQ3W/S+SoX1eC8AHHE66qle5ZW5sx5OQ3hpNFhsh4mwZ
MluI6oqH10Qd/IL0pM9R2Y8YWz01YjO5WyekgMzsEMtqbUUF5pou+W2ssssJ8G7BOBEeev2eXhWd
3ZgJ2jwcT6RCswMfgKElfZQ5IQmKghL8FZiPPXs48G0h75VFb65u6Pr7415i0t/U2iT6hInqSnAT
6rALhTTnNxf1DU7cbvJrJfJmm5cvTR/mARGVoHNJ8cK9m6WOI60AUGoDhMrT1fmiRsck+p/n9ACF
4fxtif+HCQzIse8pG7X6JeL/R5Rwc6XAHVIXyiW/Mf1RGtPyIxiFkZGnKyensChCvqaz6yC1+Dva
eYTZtnqWi2zVywrwKiFXeDeDleVqukw1ySFsF6LYP1XL8YxgXf57ISfa+waqvZL1wu/WEtCyFHEX
fCG+ZgqEwJfv/0bfbuGGbK57sjE6JOw0Sdyw41FgZl1GbJUKlvPGK//B2icjoyWGqxGSuPudTrR0
20HKyUjnF+ygMuToIaZG6+21rTkB+kpkEhvMr+opT9ICRz5JsecJecn3jxc8Y2i2yG7YiYspQ6hf
8/w4mrd6NZjysyWyiCmIvuAmJBrivN7wTfGgoStkVRD1rCH4Wyffwn8pVIOptvLXa2SKh/JFPh0r
Gp/ixDth0uH9nW04GFL3TlMDIKpbU4LYv4SuICahIi2u5ST8PEUUzp4f9CLDKac3iZNcZ4GT/sQp
ptK8cvDxdzsxpdMtRpEeC6m5cEVuyS9as3SI0s3isCE/jv9egXRGc/g4jbYK/dnK+fFNPTflcGP/
9T9/ZqL80E58puKL3eQDlXz/LnkS5GFEjPq1C08V8uscR6iw20Ue0Iz81tE5GEKmKoXi+YK85O/N
d1QhGnv9KPJfgdqeQieqAgT7oYiooTR3rxsSFH6WT4ja77zaCARgJa6oKf1mFLaY9DLiyXow9BM2
b2hgCzc3J2t7pTtefIolQ3gm1/z+D9RCEMmlkFO2BlAtpX+4R9XCiTb3iRQ04hnJmF4dYeLP0bj9
zddO025xyeYNj7eklBbYNgbsLVsrjRDLe2zE4arktSL8OtfQLhL9EWse+VpDG+VjNZET3dSI2Ccl
wuJMtJ2CfiWGeJFZ2bdfbnNTrQ51c7PVnawstTaH26x03J/q8vnlQMvRsKiTJjcBJzOzx+PViH6Y
r2SnKX1OpQXTMrQZkjqtuYZcJiyTVOScTPABobMSkQnb2FoTs127bqLAg3gOp7hybr86/x3fIhoh
SitGIap6b7hWxNHyg0scjn8jptEX6jrg5jh+AvSkYDHf4FEj5npwBWW05OEMoUJTz8TO+kG1DE7L
UMHeX/tYeSbbWOAU+SQbcpsWZvxzPtV+zaBUSXNQ8l0vZgpa5vJu8ze6tOF7no+hTrtidVw3n/qx
3TeVd5Pi8bHWNm4rAlmPSKCnmdb1qBe5cyzoomumEDJLODbSSv17GaYQKyK0o8Cpz1rNTvdyBqes
xgBHIXD0gWa/Da/d1e/ekXJeT+pA3GZUtt9458ViS2wcPZVApZ0mtKBvxxFDf3s6tE4IS4p9xXnq
nuOPEKnzIyxUPFAr5jDbozhCSpjrmBOdNMsi5tcW/xnS11PDNszjKIQYfi1h2PyMIi8eeJS2Wo11
FbjlTLiC+xPkBlFIiLrwItu5sEy+P5U+wfbE2RtoN6dKAmq9C1dYvgnFFIMAOEiEHqohvVfruPFq
halmedsQHIBYTZ9nb56swsaAm3+U7RqWXIRl070BnN5LLIlXOtBbE1cU1EohwkEhlk6qolqQH+4t
CQ3YNO1xHadwIToWCTVxF4vtWNXSt37O9GHMwtAVlm+FgQlhtRkaBvkIEmXTSSf2vX/FOhItsea4
yUsnuauWIAQZDnlg3LWO4P4StBGpg8eYrjbEggHi/73mwEezFosJLmzSyZdVBXOhHsNM+nKrdfEH
R2352QG4FzVouiuRUxWFaLLdZ6yEwreYLNB9CybpT+9IW60f/HO/b52yIQnlIvFnoEJCuvK+NThx
Weos1r//Cv6n1dbL/NHLT+f3pFZBJ5edfWBPneQsIeF8ATtBu3WV04uakOgX4XXRSkQr0mApeQCY
Xf4H+SQVIwdg4Ac8dko+wV21l+ghNl9/RbytgrI/d3bDacIBVJVwTPitwxrVTDQiSJqzTRql+92f
DNlotX/IfmEfanBi3Z8MWkXaqO8SWQZ+CcVFCDaNVQyLWy16eBGvVxoGO/3ozOZJ3d212+Ds6mya
ANbX4G6VKxpb8ctytaQDnuhWWZ7HtNCxpaXVkhZjKuJCgURW+kQhJ+Hu1J6AOffj9PFCSxFH0vj3
1/p2xgHHwUpW24lZ0Kw0wOdcoVUj7OVmW2t3kzSED8pqOHLUW4ZsmXXPm8CHImwcoDw9ae98mvi4
C3w8tRI+g4EdiJV5KrpfUFwklsGYR8Xr2i9WT/5fh1EwUuPOj+RhJO/90Cpj4rL/dMaheQ+rgcBR
7NuNQ6y+YfMuYJkFUux+WseDi92HcGYCOjwUM94MlXluIzSE7m4buSP30wRcwzXwQfGNdnuPkN7Y
/IfB1w2LBjNKbS+fr5SmX/ViquX4YFnC2m4Rs3ILXNnrMwSmByta+bBaHVJ3xev/oB/XVxrfCX1d
Y4W9Lk7hrqydN6CFSNUL6tR8l8+jMmNcf1L47Oa8z5sPP4MmKNFQrP/lLO8viULVsRH/5NQEhdAg
eEeq3pT+YV/0ZmzaHp/OlBClGlLYWSdBqiyjrlkuRr9NZSDBsOgcjW1U1CH5afbPgkFVv2VNI46u
Ao+UHKV4P/TiCWWith8am4DUIvKWYLaYXzxKym/j+rreAlV5YgpdAfi1m7jlLay7PEQUUtY0E8XT
yJO+aVTWqxZXzy8cJOQFBYBpQkd9/3Vr4yS3dVfhzynL4Qz5QgYyomB382ScaxOe+AYZsrhXN3gK
fzjJbEiawhyFr3tT6rMNu4FtI82Ohp2mdGJ/mha+LNHsjpYrC0/gKuI5qXV/+wfijGuKfSuFvynO
56bUcK7iHjqaV/fpIyT6MQPCVF5ncnksD6ChIiofY4MJXLQz02WZehpZ7mXbxhewx1Ft3kxnvCLq
FK17yQpD9iXvuwjTGtGskEj2Ugt5k/b9ju8tFiVqxeIx7QyE3gPWvT3iNtewYjKx5EuD987nb2mj
5hKMd+TTMUr5Gp1BR0rmSffVsLNwT+L7Bg5Nb0cAEB3MTgysjT37DdifUQOtmzzNc3pXxuwXXLPw
hyqgnkkZU0ffHm3xfU1ZxLQ7tyRRcomGLZDhQTirgq+ZvRyoZ8bVXETZXhHstNw4aUeFny7U8DmV
+tQmIlafdUyvVcNsw8gx1PKpZAzuvN3CayhuxpDtaDsjC5YgVx+3gCnzsAlNz8Q+xuFCux9aL6qW
37eL7pIIYCuBahYuUO6gkDm7/pNSqGvUq/iB10TOjgi8O+LyT3fXmd88giZ4Fw5wGiNlOy2ZREU6
glx+BR4Vk60DDy4PbgNEmc7yI0Trk/ICnRwG6LfvNjMxUlrTVQB1SknOW3h/6j/Z/yCRoede0heW
nLUTKnUNtPBKYfX/Qfs23cwfqG0j7omksZ6ipyb+xaX4HrpcHGZX/H3+hGkAvpd0KMILJBDT4jbs
kPnCuHnsx/jo5ZNOcSvbkSvTaVlxAWoMV7cvb1dkxnBVLg/zJzNkhnQT4C5pT0rLFHcRDiKE5jpV
Dttsi0kU2iiMveo/1gY2q2UZUEmnHwAin0msPHIzbNtfXVnk742bKdjKjT/dAHzzVbIn77AUtHC9
zXgVqKS5xnIcckU6tm+bciyZIRVhos+AlCMI2DJaiLkcoi7Zw0Y9ve7bc8meLkfmK43rVFZ3R4oH
q17RtntZywzXktCuRzMu1GtNsahUXA/kywm79YiEN6LZMNmYvUgDPnBy1i64Y/fxYB4ydP7G5iRe
SIZUloW91SdzVlgAOeGhLcfHef7ZnE0Gk33jz5orJd6j5YOKVp2vgGCrhFSYw2EdEKScAgVnecNx
WAxQnM1Ff/uFoxm8/HbhBYjBTdnlzuEPRkGXREzyEgO7nMlNSxaDwzmVlDmwuifGTb9Q25bxxZFC
U3kS36DsPP/ITWKleb2rbp/NWVC+7QXJY65erjQRsz9T5JVDXq6khKcyPuGdc3wfMUEBXArjff5p
urKDG9T9gN79OMlmDVnyA/W2tIIdukILjO/jGTsDD3oWODO98oGkDm1GMfTDHQnLsC3jD+Fe+J40
SKo3EIY7dgqAAulxH4TavpXe/i5bJQMXFUz8fizUeutxdDGhtt/iDWm/Q2AIz/QrHxODNSETj1Am
khMiPk+a6/NCOpO4zSHnye0QrWuN0AXu0UJR23LYjI+zfCLNp9N/vAUecUH76zu/T3lNr08laZZD
K6BfN7KNoWnN/0wLG3N9tMPw9BW3T9qFseCBValsyBYHPHqUezfI91Mex98lRZqMzwcsKi3x3f5V
bogfK/nm2VwAfmrZ17aQpAeN0nRc2eEUt3T2qPJnjoBtPdGiRpipBkEVPAQB/SK8wTsLL6+CLTHS
amPIx/n9TwhMBSqomFoAArZojGpuKNSxr6qyp7pGXl0WLW9rZnRNzsUFVCcVYWrYLjJsN8GEpias
g3CrSS2P0TyfhlwvVi9ICJeoB7o6Tk3VEOKXlx5zGxBRrIMsZvuXuCslYCOfRRdp2Bg3Rzak2DD2
IVXkETDaR7n6E+X4gZEOD7Py8bvjVEswRzlbFCLOpL4BAPpv7vjtPy9UJu8MV48okE1fZK//1hwg
RV7cyBjFYwsYQ13liT9H5L6xqHU3MtH1mo8/zsyWtzEaRbqb6OK+Vds1PIMPb5G6K1Bq0RfuFXCk
V/SvHWTSO9gatI8nTUOUQsgMJtJSKuuKuvh/hA43huLBHMkCtHJw0GSe3093Q7QI2EvkRAGGGtOt
WY3wZX1x4C/MbFe4zRZXtOmkmhgCGzbuG900Tjmjl30yGJ3PtGL++11y7HAaSuQaxLYbu7cDitss
Kuf3pMvOQSVNcrQjmVupfdXHlTIWI/5r+vL0dDiDTth/RFuoAW88R5B2Az/oBH+zGqXbXrpbvI+0
NIbwVMqCgpvhjZ2ysRTwpPu/wZQLzcX6hsLHfIBVO0dVz1kysF2XjmotIDO0Z9aPNri+oRPnV9DH
62yXZ3EG5k/+LanKz1zYCK5XgTo1eBrM/WMikb1orEoAVFns8vsoh7piss62eVf5rJTzVfn2rpJV
m7UtKecrRC9Kg4PoU456oIXJNyPhA828UdQ8MQccTEhYS+k8S1sJEL9VFW3di4XOSETS1jrAEbr1
IjV6hXPn+IL9knL2CBBRPRbbFdCv3pvNYQyWCqIRmced/HMm1NBUNzwBGqO6W2tvp0kZGYh1BwUO
3YnToirbKb1WqmknlmGpZLO1s0dP3czd0HT+kloHOamI7J8j0zVJN8V+rwa5Qw8EFEMXhPW0srR4
d79TXUPUmZ2NIlnUTUpl3IiSCg8p2gMSUblvRzfBQqG6/YeeSXDnHGR0c4C/6dQsdE93LfNlw9j2
9nujrupo4hfeYuVmh//X1SA/p04i8cZtxsoB7DyZAA9wINr6mhFxCr36MNQKGBEEfxTDEcck2KeR
iUBWRUqEdNgpimQnJHc/0deMB8Md7eZURy+sbbSSiu7vXvDUAA6oLt9WsBegnfrjajjQzya+tR9n
Gak591EmJ6HP0H/fvvlIeej+9S9HAFtmiDky/DV8TmNlNTuDFRaatV00UDtefnS4sj2B659WDIcU
Sv0kftD4o+XfliraRxyA1kCnluAcwTIMZ6VqHkz9o/sjOWk6qAOoal481mG9HsCJBvSaI6ipvCpO
iF37ytUXmDEku1XuaLGAiSUvIJ20cAKgvQQHLbotYXjpEtbgUqyFXX1FFCbQ02cAekzYYfiAtNCd
1Yop82RE2T1a7TBH3cJLKue58yFEsLaraKZrpW5kY9DqzheEQjOAhW/qdweX6tj8PNTcTRA0qWrq
DQ9KOyqB1Qdp4XJ/ZgRtg5pCMzBpoEyMTq5KWMdHb8nOXFXXbhFBxyO3R1Pr5v8TBj5vuuXu5BTE
3F38Bnfm18xGrjL8j+K2yqjONnvCE+Th5GuJKgFxYBgWSMFs+zcC2EeWvwV/03NVvHFbFSzPmecS
RahgOM0I6saviHPczsCDSUpDgl/nX6ZKnsh9NaoefWyYSORQUDJjDf1sBs4nabuUa3/rDRoW0mbT
J7xc/C12i+h+OD0B91G+I8P3CjciwjbYZUtUSRRgK0trtohThvULO5gozmlQCJXFL6lBqQ+/8s9e
e1nrknyx2mGPXdDhMSRg1kcTWdqNwIOOe9cLNpsmgk5l/gY4Xz71qj/LB9VAYyNCHoI7x3LtEq0z
BbMm2NzElhsgZH26wRDoqtV+TLrapmrrIPR1IdS+Ev1u4QztvtZM8xpzUn/Sbdy0Gc2FD8hY8cqs
cvNmOyXpPhh4P+6V80SAQPGroV2CEED1NOEBmQldf5H5IkRikTvGY7GDRsCHZCKb44sYuTYL78CB
7smMd5feb49RiVhfeXRSQsFqwbge64XJykFbTwPWC2MkP2CJNgyuK0Lu1OgCIDFuxiNkOtv4IMVH
e/6+H1SNQFMuau0H0LGZ6Swadsuzz8Yp0vTJKaUeYjmDJA1dojPkY4+vRDRUXZM1hMeLFqcD4Ok2
dKThWxUXaTbVNPiHxq1KV4vwMp1ayyJlu+GozfOJcN0+JUlCNYRbQdYNyM4jXaMGCAWXDCrKr0w5
W2IRjUChnk7MDArQ/Y95c3pIxOynEMuhXAA/dCs6HWk8q+/BUNefaH2sAhrQQOziHw2d2Ia0feNg
9E6tgUzylCmaE39mW0b8BUbnY0Cw+0tmdvXuGNF2DnoeaHz3xqRVw8dbxuhv7Nq6V5iKclaJAw4v
OIem212bmDxGn6g2mWxZ7q5v6nwMp1F5+Zlvts2zImkqiCjyO4Cp0hgM/aMDAsSxSERKJZDk0yZs
A6rreUeGl92UjeyOsyKZeABZjTx0CVsK3+RU7+ZDY4XdDYm6tDnLvG9ecoZ2kQ6RTvlZ4MbXpyNn
cAbqbaD0D35tKO7ScIF8LDiGdCHsTMcbiqQe2YSHzvNbRQW1lqQryCPsQpaEfEXN5/x2LxtKz8J2
uwJJvlwCV3LvXk7CCRHi5UaZMAUfkMWowH/KoPH/n76fquyHQPWeWxCfZoInuw2PIdPEeUlrPPgP
xBQUP4yTfbykbKIx5vhnSGEQghEHPuCdfR88qYUs/j4N0fUFaX5NR8xehmQwxcpwqafaSC7osYI4
R6dJPSwIsoDGF3HjWAn2hLSqbGat3y9puNeuCRIc59erDttCZttd88XgAO/el44qtwqHlJ7s3U/J
sIVY1RSRIp5uq0Aoj+DzUxhabmWRBeIvy0z55fUZLtG7j7e9evSd/yRXA0DCb/4ouHM5QJjoySqo
5heOQ9AKxG5V73Ez15IHi2xeeUgoO1k6rZ726y64iPEhWyOFT9UIEHYmfQApaRorv9PPqpcmBv3P
F25qUjaIH1PBqNtqYkqEuERC00i5Qiz/3DIVsPptqsuScI7qiapSAFX3qmc8JBSrshKjgtYwdUMd
v6JUUbTRuSXrop4Yd62slfc0aH1tJvXIqzQJCMz0C6eTmQDelzaa0Idl7cyk+QRM4twZtocvb0zT
8utdNvkr88zuqtNa+u9tp7P7z7DQn5OWk+JAxRu6+zcZZ8pVDjQSoZawJTHDTJOodmT6VwbCjkdV
3pIE5KJDJ56LOVtLXphZ5dFqjVDyQssfuCzwGB00UHwvz37iHgAyGIsYsO+JOhWDWcq8KWYdV9s0
uLmNVkMLoI6i8RfrtpAZ0EikS7HS9NV5xLNh9nq20lFOw/Lh+75OfSwPcHqdJrXrQKQ3fZ3tuVHP
Wc5vSpdSMdjJ1OtDwHeAUfHs3zo4qKXl5CLcRYVtgjjYBkYVh2vMMsJfFzotFgaNWUhjI+CbHbh5
FduwjXwrSXgxvqALKzgAb34TzPvtLksPWs7imc+5Vs1GPgtfU/go0jC9UPdED+wfrg4Tojk7HFsP
ZqRCJlEGQEBal0VyIPSDS+6ggRgFuH+5i3Zz0Y+iDey+Lk/91GIjUM7kUcbipL6guYnNp40I1St0
PxogHAh7kQFannoV/CJyy3sbqYwDIU8xSk0Nby02MHlbz8qYbaMHUWho1yO19U/XbN9ONFSMLR9b
M6hXDp0PXpXwKd028XYgak/ETAw3VTXmlV31Nw+KbEIK+UiF6/UWSnCBgqNOUlFOWuRf8azWKHsl
Z+shHoBhAA1LHvJc8dfvbbl35HFNWHNiNI6kFF5Zla6v74ISGhuypGMGZNbw6lQRv82g5VUYLoBT
SjdIuSdzoU42de7B4+Gf2JjysGwefnk4TOmjrUrKmag9ZwfMnKTLUXu8bJM128DGDW8xufMozdKS
ICj3gBy9ervGOHr6XdPOJOjHBGqEfXum6nScaX4zEZ01ib5EomN+fg54YXXhV9rPWKgpPV+yTT6Y
5kqSle+U10sybAi/qX2UQ7wPr5YRZbRbcVCkVPZBxasqY8oU4EqnS7edzlgvQWkXgoOz6pQhJJWj
xlzaIDp8ceH6BONR6DXBWzRmbvmSpwyKKmQ3XrBVM2KPMzoQCanKRT1y0XmaZM4EbX6aKRlD5JEa
IsXhW6Ef+6DLWIHMNJO9wEFxdffNckJBeVNVC9LSm4hk16uOvZx8zrtIzo4Dm2xi8mafP6sAJ1QC
8WYdhzDDF9Qs8XovRMgV0faBlw5eYqPArYfrbqC6kNnFrzCD/hYZgMAVsJWOZx73jJrNvAKvzkBt
hcoF8fnHWI6uN1UhZ/TTjeifty3ChVbRt0IGGdwdO5xMA2NKVJMcwtpv3UlODmoIM67mUFPq7xkn
mFCs0cB0BsUzRpy8zx7T2z9lWNrwJeNc0NGsPSVFbf7siBM+mBKuiz4AOaFi3k4LZPwc/uXoLw7h
4R0Q2u9fxvylCYgvGhLJBfvS5HmYPLvjDmB/kvngXiQ8Q3yMjEztfIz37kHuEQVfMXagnxaMzjw0
KSM9EpuUo9w65325dZsSTUBrBsOM9aBe9oyH2ZXPKkVmqLrOm/+EBxBoTRP8BlwWGQfeSqtGeKRl
dVcOz8UJrD+UbjZIigK5QLawvWvF7yHUCyJy8Dz8xKV59BUYlAEqzoC5sz4p1MzA1B1S2AswSEen
kPuIj3UCVT6QQHCWmTzpvYc5AptNCNYzjptrj+WWeae9bcHuIkS7rvex6UFf1wH+/p2TGOitWnOL
mIhNDpqOgUpmc2Z1CkRwgJzx2QIz0M4310FOCs/QkZN0RWMQrfsOC/saYrwR1qDpPTdOz+2eR1M1
KAO/WD9u8GvwdE6khqg7BsOQKOgDzG4lWY7H58ke9JWpgfwv6BZ6FnughlCbwd70FtVhbUb/7x8J
dSBI/kYNZfcT11hmc86JD6Mtf9twM6pcIydDr21e1nbdL2zh0T/lB98fCLRabQvcXX8mlptbRwch
qoKK91Po8TGM/hKtwAwyVYG/1PdLCJ15WquStch0BaKULVctWMNf8y7n7NpE5M9PrsK1n/TzVG71
qnJhJFCgD1VW+wEtLZoWAkPnPS918v0fXEzcOFQj1+PkCtd4Dgdje2V/PvGl90NkYTuHHp4pwlDA
778z30zuK1fq4BiVIrl8DsO7P8rrSflwyPBwFkXJaN4AGeuhxlivg8A6yandtoIr5ntHN8YQEiZB
rSEnGxile5u3+21cZapmptykS05GXU7I4RMexYlt55B97UDQaEBa7n3p1SawAjKEsCT7Gc9NHwBB
OC0CGyJ5UVpc8y7GMlN3Ia0F02tW5oWGJyc9DukUwGo1ML7ALM3gtmxqbaTmNZ5a50Gp93gOkSFj
vAKaoY6+TYscNzDV28GDUO4VAJrZieqU+JBLPRaTURzvaZ9mC3b48Zg8lD2XtzMeLXK2xL1AKYwe
0ZTu8sWK2Da9VYOhX5Z5feXwQocoLKWveECMG2Au04mRgD/HAe5NVmtX3YhTVxiwe8pyDzY9bvPr
6xN+2qSsGJ16IzUp6P8HGbfxaw3DLR+/oKk/Xp1ysoxCxI5NRrNb91L1SnPyy6Wprk/5tGzT6xUL
E1zOM+m2D8H/YwzisUUIAASdr77HgeeQ1Aoj2aSFpm0mOriT142EZkwXzKfD+PY+vCvCvuhvfP+r
obk6aSuyvQjskofKgeDMZkwFauQaSwg4hjrV+tJYOx/LeCWDQDFFNmYzbPLmC9w6MlnsUrB9l6ng
rA3RMogxd71O3MaiKFCa+lhpEgiCsvUxuoQoKxKNNkaPTI1RGGzbdXf/t0wP6zCmnEvqcN1sYibb
0NNN8da2Ramq+LkPTt3czItOsrqhXcDg4bGfHnZWNqViwRLBa6a2DtvpRwrLhfv06Bxesq8t+gXk
vWsjelYpz3PCg2M/oPuX/hWk3wgR2+tf25/5JwyKMKgkqlOkb93uxRO+WKsTj7NInMj8oaxFu1sX
7FmmN1km00v57gpbvnspOzdzXMAD+045UHNQ+8YkksKb25jU7dm4Eqs9QLs6xfjPrhzez/Iff+9M
6wqOB7Qbe2M1J9G/HCXanmPchWxA+FBtpThI9ZJcBqBWAA6JC9+qnVTq4kZLVhxIYBcQNMMQDmDN
vQ415EyRU0LyKgWWDE7MrfQPdC6aMjp6984sEuI9RHsfxUvvb0s4Jwz76lu4wNDvNAkELuzmDPzw
PBdDinYfXIofFN/vSO/2IrLjjHJZILIZGCmxH5PpgqeN1rlVbmfZMGvS8FzOcWxGY6cM4wDZewH/
O6r+a2yD6E6CReBESCsYw9Q4LapvzhTA5c/ci7DwVxdbvPFZ8RJn+wj4tVYgmVeh9mMmb5gCT34P
CWMaVC4nf+e7xonpEPMX1rOFYyAS7TAoCAbmyvaMwv6d1NKHvWDKi55WIFHCzREfl19Aohag7Vf7
fpW7uAxVgB1l675up6GmaGQi5AOSn2vZ7Aqyb99qFUF65G5DZBFYyz9s55Z0pfrXr3lUZBcFOaA6
sLB4G11pHovn+g88zNyFMKnOiNGtiKuVQkOFuekWwIhwnmlSOWb7Kr7PVKgcD3bCFl2+RHd1/iK6
wisrjjiimsIzpHREyWbMC7l+99Qgc7Nm9PpHzofHiX76GkqY4Za7xn4Wntz/YulBrU/4WSqin1vI
JKnMXrkie0+mzrIvY/UAdlWkEjuHyTS/x/JpPIxvnZwelUmC1MU9nU34Z+l504MFYpG5IpTIU68y
/+HMNnY2wNXeljlb4FS8ZuDpDqn2vZsYh/LgO0I6Yhd7VrZpSr2PAnokRJCpytQAchDtfHA/ocY3
i1uwlUDowEPn0wc89SC09YM1V+kA0T2iacytDci85F6u2G6lh7wgLG1zRRrydppU0ND7SFXvdQDF
p7yoqd/yoscqv8tq/NhxH+e5MCuDQpHzJVje8uAc6+DKhuqTud6qRdW97zN0KibEHzvqrhrK74Rl
ydzQw8zlJFr5Q301mNsKRFkz4WPx87IrnS1QlCPNBC7y1qsF1SS70Vqkd0Ft/XCOBFyjeSs6ibYk
vGDfJwpDK4RZv2yHYwxKZH2HuzJg151PR2qgYbOIbMs63kM82+cT7vZwg8/c2z9QN729t+B1fCRB
HIN8HKOKENYS47/8W7pnoQ6mghOFXyRv4MvqHal4uSeEBOLt2P5A/AuWpUe0IalFGZ3FhNkXXq9t
coIDJKGL+8SHk4W2jCOGETHcLr9twF7ZwLdWJojWvJYtFpI4/c6tExMKkfxP+dl9KGA3KqF/3RWf
DaRjo9N7RKgDhMLuULbVgvn9EASgSMLkk9l0CBD9hPMB40fWk4IOAVOOOIccK2nhrDSst4Pf+Jm6
P8WOd2X0OCqrlQG6jCjeN64qwzrekEdbkKJOkeMLYu7Lkyw2qcrBDB/mHTSAuER+N2pyDIxMq35s
gJLySRjw0D9ojJ3HynJ9JyjDQ/dummuZUp02mq1wdjbrnrQ/lvhPwTVVGNEwFGkLkw2smANkRLGF
g+Otn2e1X9ijWEbzVoUy6HwmZYQtsgvZzXUGnZzJi1Sf1Q18RF+Uogi+15qda2t3jAuyCWp2ORhS
TuPys0iSO76GQQAaKInpnV8dm57Uifbvm4pr6n9wTNMscPPtdMG75gaCgi+wsocKzIIyykxu0gk+
GroSOAbQmxJHizReP3lYBN9P4u57nphw2J1zKIXzPUwUoSrvN7rmG8fnaB8V8uMNl9RaMIJmY8Qr
OMcAB0coKKl33DLYBm5elA3bS/YZl/sTfySSdcYzR0eojpjj29NVh1EGmOgmMPwEBwVwL7dbNPMT
TBvADgImWj3ZW4GAORPc7GtiUbp3FOJnEwE2+/4jOb8z1JZq0nHffyyrUAtsAz5TtgxRRpq/+PS4
JE5df8atXp2EH9Ddor9nTZxM9UxiwcdObB2m2cgCZ5ujm5q6uJLhLEjx5EpEnCOTuS9+OSOCvb1p
/NrEcWAvDatRYWijyOitkthMWykyAe/SEKYoJIhTS3OW/pIFemL8BMD+IHoxb6ZZZl3pN7J07UI6
Oymqc3yzmoOP0qK7E8LvLeaefqN/myADDVAFGHF8ul1UoHWbaXnDl4oiCdeBS852x069ttX61Gjv
4CzBcwGABk9Ttq25jMrVy+34BVd548vtK5oHurRzUgvBbNQSjeBZTznmbmZHC6TkeVBzNHEVJvb7
ksVUtaMoVb/wOV28RfxHiXWaK51drkjoaQDnIZ66gbTpBCAWjqZM2gCYytWrV0Bm1XhqmBXYzF3h
a251cJPN6mq9FPfSwYBOPB7Ijjyqn46jVAp0cnphbqTqZH9e/ByHPhyxE2msVzyvLaFEmnNJ3UI0
ooHIPIpZz7XMp6m8RcykhzSwbNRX78i1NvWINYKCH+2SaGcefjx82+V4D233tREgVDJd8uupoq8c
l3u+2rtF8UV8SWXoTd8IPYXzJiBdiM4KW0zQXBe79FM0Aba1k2TP7WQN8zLesAl4TgzbeCP8SLRC
V9Mn5TTDuKgmtQngEKN8IVe4NEPoZizreQP98VcdGovkjoeMonF81lCnyD5wYTismZMTpDb5b+31
tIuCKbGGRzvwJSZ0dlwbCxl8Fymnpja9PN3FeuVyZHzjqv+b3Jr8ELqUy8biwrrWmAXuSbvfUoiy
64lE65vFlnxEC4XNwFcb+l6UmNTT+q2fazR9+TP0Rjiwa4cyMq9FBoGN0UltGQFq2r7Pv4Cj6BDh
DR4gjjbDzkBisiophjqLSecqXPBFd910zVt1Xsfdpexp8j1+F4D48GLn302J5kdc0sITdN5YG45C
h3veHwpKugfcMKbmtcEtvWYuPzFToBCSlQnJtRumgz0pfeto9Z8YE/szsf4+vWUW9J7lbhZLsji2
xgketkCM18PPSQ9f1vgpPSHjWw+BP8rdX9fbavm+yGXstIZel53HZ9G9U1xzs99nbCDejZdjGIU8
WtxHc3KsOqEgl+X2pQxps3ZdKd5AhtA5PLhjtGv6Q7Tn+0nGyklPHlKFIbkK7F2TmJNCvcQxzRJ8
TAlTONcL+g/b+Noqk2hjJvwqFEXY0uWnKoIhrGqu+4plch02pv2IZjAWMWz4rCI3qy+W8kpk08iE
fj1HZR0FgVweUJJHuVyIqpbp5Q7zWH+PENlOl6PKI7QxufMqBt2aX0wO6LL/t2084eM4tNOv8W8Y
o85oT3xwUbX+w9y2dXXPNDHewdu2jWsQR+WhWs5CGCILX+Q7pHWezUENQEm5QOUsXFgHa5ogFNxa
1zCId9sj0RQ4wJvMBAIUAkKL8X7U+Io0bY43tsCN7+dL4OSp4JzFruVagxhfqU+S8whYJpmandP9
iyEr3mrGeiRJD5djk69B7zyUKRt3UnEbmIfEbzI4P/fmEFEZ7NqYjzIXHvaOr4l45+a3GHJNLr5M
baUYcDTPe9ufAPrrlOCQXiS8hhO2USwS+Sxp3q4thzoT1byfgc4XxIHj7QFVfkHWlCIlGKNSbAp5
v2lkTHjJ+8uDXm4cjJtDFChT7Nc9TDJunTDgCyXOxg7lyAUihBT+tAGqLkwfWnTPcTMjOqfKnWzk
RL4Gz/zroNW3Uh73v2L3eIkDzqLeg6Xi4UnFjYF3pK3wuKFIO//FznUnCdZlBd7M57JYM7h3B22Q
p++mSk4k85LwUGctJNgGTED0mKHCk7oUAe5JtinBcN21dAST+RKL6WIWc9eYKPuwRKUL3VCt1Ok8
IQdxxjySajg/ooynjTTy/bmsUQuewXnUKI2BPGGfK7C+A2SPJ8FDBVO9qxmwfBJy8oDZsV/Jx2qT
hXHkJ5JeIDo46wdWQCwU8X8ZZHrn1Q8qoH5rO11/DzMbtv5hhTdEDpMcQ/vheIsCC5nYp24UK7qP
O3+Y1dSR6sIG+Y5ujBAcrmkojCY3qGmbH45ejXV9UT/xV/GUZzaQGsAGtSza7AGpJXJ9eicpswwF
9pHdaj6jUq2Hl1row3Jlxbgi0ehrayE8q98s967aa4jsSuBxW9x7mOqy4Lwd0P9WodnDljWL4dcM
YudNuI5jGFOANjnBUrxYtBiUoDFJPDiT8xTpYWIAdaQA2HQKDgkWIeCH2vzIpxOlEq1j6Fk9iA8Z
RzK6tT7oVCs88WmfZ/Z1W7aflp+dYwYp0beaj/zNiE5ktKLqm9kHRaqsBxRUMG9oCJMm4rdcrean
xViK/xfErfT2F/TeodZhW4Lxpqu8h3cO2fwngd1JVFQLawe28zqQW0FXHB0XxxeSvEVulpHCXVcm
gOkuPWpd+Juv5IM7fT/ccJqzo01j5nukqVZqwIxfggpluVP2Cxs37l7TXU846rS5tUe31ISY/Jg8
N4NOVAwtQgasbI6Qufh6nH8hPkd8QoYHEEs9yT4bV0hlqvJsgdMU6VZwNoSIwD1EdNevF8hqLfTH
JjmK2qdJijKN+33spm1xwFCGFleu66ckJN4jCGUXjTaXXCH4ySQKe04IbgnCs9NrFqJVBG0Urtuh
SGq2MX+1pyFMTOu0bq8Bh0J+EuyveScRVkyzO0kRjWwBWo8TfTBfc6RJRK9oAGILo+iGxpnURf6d
cOb8heIEEo6DcKyUUt91pw746w8/f3SysgfCV3346gOdPJkSsAWF/gL63UdVx4DsELzUbQ/3kut5
8bsCzoLPAz2GMNg438bNNaWYS+mpiGPL7qQ8lLU2YDfYgRbvQhoWpPJnsNlvagWMdqT7V6Hagbuu
wai1mvAm3RkYv4RSzeq1xzmAJziCrqDdE1kz96kwvPlSpCIZhIzv1xcprOAKxT8LfHqcvNmf+L7y
piUAHRhaAm0I3OkOaxZI85dcanXHF7g39yBgA55rlPvyYiQFn2xKsoWFcEzM4ykbucevy1rA5GFE
xfoWobGr3/54kOiB9pWm9lr69bBp66K8Gj3yZoov9SoRKzMzRUfC03a0ECJgp4WZp6S+Y5VjLm/5
k1vDy1hh4WIoA/VGc2Lcz14wHErOToe9K+XPOvgazaBsNqbMEU7JW2d/2l8ojgZZlQ7XWCIgS56z
uoifuGWmqp9fsL0Qa1apxWYbpJrytYmGl225+nE3obOQ5NbquPg22uTgZGRs+0sWARnEVncsyeV2
bOYNMFa9M3GijVDSNWAffxSvVY+j3NFeHd77nTNE5Y2snHrMaq8dz7GbsyjJyKcQkZxO3seHYEsY
fJxqWJ7JaJZgDqhGraeTdtirgRo5K83Dw9IwIez/heQHtiCGSqvkLLTnOEqFsNg/+MSTxQF1FFpf
7EE4ZbRj0j+bdIYBJ0OhwbJFQTFFjX5oJFYhn7Ispw3Dvz0kSxqja5F/m679h5k9vQ8u/lItRzbn
dD3u0099rk2LEbHX0NE7PqX6dwm1IzBtkazmyM8pbSjmsc9LVU/FRDnWHWBLDbJ4ChNMJf/T3nlE
FSd3AHVDJkLRWPvdHpWDaZkZ7KO5IMsnQmmEy+wic0HpEriAG5UPbhfKmL2eqjrcA9KFlxsPiwLZ
UvB0BuBNaZfeh/XHoFAuA3PXsscLVWS/9AHT7rAYbW7Er0iNYjE8cjzyO1Kl0qWBE1aFGafSlnmT
IksKffQmkdarXq30d9POJSpPW8MXD7plpWio/hxIxPs0xu7EDv+PSP4CTApEvJ5eAGbunnYYeb2B
9U8x8xoOs9p0pUakxCEKfBJheDUnhlvmh6BMF2tqT0KgwAythXqK0clgBgOYJQXmXjMUYTygZtM0
MV/QSFF6OGH1Sw8wXgffjr0/GskOB5YNtOH2b0PAnZtW7fPFEeoek87FTr3koy+d+Bel99oG/zlG
fg7s7NDyaAsEemBzDvVeGnTlwW4QZZaiN6FG/we1k+/E9AGxNyFLGgsUA2KCpuN22htE8O2j/0nb
8zJPeE2BOmT2Lyjx8aSklauMlAxNxCbo1fjBabBlY9WKNNIqW3vgmgMpV9/BpNRW7ToTkDfF2bBn
ge2SVJT0kxSxPhDjUi8Y63eAkOF+YwpNQ568fXu8nPPjvJRmCpdVlv0dcLNJS4ITyi0r8fdF3B/P
uuNnl6EZfTgYrMrj/8fZrzSdaWywO9oGTuHmlorLNFjH6wtTPNcuuex9GZqJ8BvbLGag3/rATXzH
cfPZkO/Up1AyvOD/Z7t5rIJxEgZfq4Atvfik2bAkg2erP9OLZSLNq99QdZ3S+L4m7ktOWXiGXDI1
JOnaPtV9FRQs4tnkyopqlY+0G0tabczxowjemuF7RgYIye6SziXZBo+9Slt0pIiK3OBMOlUaVSS7
ZtmVNgUr+IYiMOHo/jOaiTFM7VYfrzIcDeE2gaCWsbSMDGy7BwwQyo/XjV8aeD/ZWIybA/MbviAm
Izf38Qx2lxPOTv2+j39be2Vv/sm8rV9OZjmQeWrn0B1R7OYBjnDOl1c5opliLIF5wJQ2G1ZZ8aVP
vu4ywTDbR7aX4ph4+J6/uomGM7VhupVeMaA+PrytY4CHpSf5QdqVsKx19RqIqpOd9cpmeYoTz1gR
efJkD3fH5C5q9CdttAAEosdLjBkwAfzBHRz1WRIqV/mwum6tWCcw16JATdLgPJoNzgHzHAX7LlUI
myWO9Y8yMmAjLxTBGDYLYX8IPeW0sj9lMbpL1N7W0q6oRqzu9L9ZDkQlZSmvSHHuC/6pMfWeQqyc
mcpqOnMMfFL+sBapLBVgzJX86FXxgZBqSmF/unmj2DmQYoXAvR5HRd8N8dI3FdX5AVBbOMNsszan
uehiJmRUawbkmNS8J8z9BQA11w/YUJwzdtzQwQ3axZHC9RZlVAsfMm7POH/AMA1muQ818prWnlnX
xcU9hS6gy5o+C5EzMQvBfo81Y4xy1PY7ZNNWRelNuL0OBo5KTlHmeQBSNIGo4XQCxs9CAEXTlG5z
nv1CvaEtwAbG+WPrc1rvLPzp1ehIznwHejWyjtv2uJpcUAIhcgLKxz5irolmSsr1+oPBrWFE9TMk
DQIm2qkOIXQ8XEUPmNPyPukATSFV0z3LAx5ymIW4Y1C2RjsC6U8KXky1VmVWCMhOhD12Kw84IzR7
QNyhBZc9l5wQU9VccUQLZKWb5CxYNZ3+xXN9s4DCHV99RjKx1gE5cOmpr7xXo4eFO9VsPk+Xv41/
/PzP4EeMG/bWjappNaHVMNVB4uHw9DtrCQXyV8Px5nHll8GFgyu1G0K8bLIOlDnzpPSQhYLNmQGv
VdHPLW4yDnx+SQYpWMTgW/uHHAF4B8dPGSP9dP5W92yf9Nkade7Byy2u4vn/t7vQR81o56lOhKa8
/+7fE7jE8Lk32XXbdc6k7+gnK0Y57TjctVKk0M7+hFnltwwp6+cnAfV/yoVwHGZojtYKhVuH+sfM
bCw2g6pvSOy5GOBjDvcIjXGYf/04nez+oO6j79jJTtjh469FlgQnhsdPuOhI56KIVHETp+MNd7S8
yUukc2fTsIwTPPsdFcDCcBTBeQfImjQi9qxHZppzl/ncjaSDLVQPaGKWeVSf/9dWw8ZM5vJa0kcQ
uRzgmKFVwJhMa+Fx79fB0kOka5ElcHUrp+mJ9u1kOJoRz9Y84Ymwb0412dihKZxE8PBsydqMu8lk
gTg2HBkiDtfSFhtka1fYx7ZwcOnUS+aU/2bKXv7MG2XMX2fL6uu9kF1y0gwgzX+H/oYfJQ1TB+jL
LB56MXBVNNIF4iM+hZ9ttbFjL57wJ3lDYbUoflmc0UxErCLdwWhQ7v9nMM8lLszSNJjqGQGKAXX1
efF8dZANumDLQ9H5eCpWZgVGOUe+mHGarLE25rqXMcc/zKUqBMIYsGNB/TFEh5z+si0tPhgIq+G+
A69omqVJFJezyst3RwjRrhNedOU/QGqVSZe4rkaIZRCrhRP952Fp4Gx+4NnGUNzIVh1Fg7i9Y6Ae
q3WjxST9LyC5M3GjAKHP+XBIsLg9/Q/PopBz5RNynMgSDcTeYHEnRrIeMk+fiqbR80ZDO2roTzD2
BRKYxlohKQvs/5pkNv6Gr0Gvc3ywIZ24JGBWTOVqEh0im1Mjt7bS0gUi0krMOZnxSASpmrFs8qZ3
gVZ7PDxtgivR2EtRgAT5vN5Iv0dqX7KkfAXYnrmRvY7ZDsd+t4O7iAtjAoOhRQ5+q4iQwvaWb+7z
Axv7HYm2MO8c/QEp/Qo+W1ywpNGwyq9NqT5YGZyBgtiqLiZo7QxnIAIPGry28rdBd14gXjjxRq5N
9EsSUjdjK7xAZCzzZG8y82PAyrp0459e0+dUvMYQKIJFEKgUz0IO/hbmVgqnTJA5W3w07GXVNb93
aYS9B/4C95g2EoBYiaIQwMDeTcM3qtiUM+64NB8c0zNxnZRYHVk0kFfM1pXw7oVMVzYHarlUuFVV
dLu+thVo66MFeyO92hD5TRPl29UxSaclfVSIRDOWyasjvxUMN1XNdIbOjrPxJpHRw4ArdcY8WMxJ
CuwesdiJH0sEi5SoeJxIMitleknl/l9ZOVFLBsbZY0miXKN3dT63dh0EbuUe1NaFTzuzChmeyLq0
q6rF5lJ2Xxw7EWIKM/mlzz/OzrwYZwWrvLFfKLgjCsYTHJi6rnNFsvKBDRVGzu6c0CpYu7eB3V0T
W6K9Vr9X4CLPGty/8pUeMagCuzz5bviZq2DjSRI5b8W7bjrkd2jSFocZUUuDs88DqrznwpeqWeu7
7EUdqlZ8tA+bxqBQu36/GWZlkrnlfOBEF9UeitpmNgOwIv0o8F42TYYHTWV2rYEQrN1YtpQ8bKas
RztH8sxKttTks2n+dF5oEp4jR6eujACLctiXa4iqkBV4sK+ZOQayaGWPhCp+DHHBS/y0rFRd1qgi
90SN6xBPrDTOwgRa+rtMjYLUrAB8oato4qpC4cQLbuNbXPqi5q9JeXLc/dNf5pV1N4KPwqxe8nVf
4bJg+MDeWnK0F5WTJ2w2PmriVFRlvHqPGTMQKg4/UeOjEMqOcVAhv8zc+0nqw7fjEBhq1yUFQFz/
rIlNGygerJfCf2crOR7xRZc00v3KekooUsCyk7SWNg7axKX1V01kZdfRd4c725yB0fWwrJh23OLS
jnGPnvJP8/qsTbmZLm7FXUrE0gK8eVS1N+YHLn1GKZVh/xuXwKb0Pyr1ud698YpKZGKBBdj9PquH
iIl8S8n3LeWCX+0ESeF+qZEwasMLNYlQe1xOjH8+sXnRaEK5aAnGh6E1yY//II9ZY+cBcDmbFZ9W
0cH+1GIGLoUR8rXI3ONyAxNfVIza5WbhYhw2pRZPhEr33/9sTK0vS6/QRzdPx4I+bHfT8qlX5qUQ
AWy7BcUBUYUBMJk9UjcEziEIe9aTQ9aZVd4QCwKg4vDcNgkm+2zta1Xui/SbzHUPJgPobUFlGdmN
gb8vetpycPnKhfItbUGAuJTKFAT4sDB9NcwvzWdVx0Rm0aZurNTlUceS4HxooMeE5QvV7TKfEwNf
ADUiinfAZjv/qtW0ZC2I+TEBu4YmXo6Mi4S3KZa8sS7HCLoXsODWtv0CT0OjLrfLExYuRxNd1TVe
f24UMEzx2jHd+ayESVf+IU2RUG+mSIeccSL5JAMCBuTHgm26d2Bd2SQPgwqEulcqG1qq9/0BiyGm
hStPkMGqenP22k3wzgpJUgqknaM4Z9IDgk+Se2oMhG1Fqmq/Vcp5WxmJtUlJbiwYH9kAl4Ih6/nI
XutC9wV6/sr38tBm7Mb+ujWjAYXmXnDX8FyHd2aTlGW44wvIoSK/rlB/X4uTJDhRetFEwv6sVKgB
TUdJ0OE587w4XX2U4lVztHVqtZCBRYDi4jaANIQrDGd9b1d/5m7b9wLA8kFaf2k8Dcqd0XAsOjjK
7V70/HfNDp3CHdS9A1SS2IL1yeH88ONZZQOz/y11nwdrvbYI+NcpYCtotdKHI9FFhvpIFMw8gjXD
B7ymE0al0Golk7uOHGUaiFzGprHyCpLFtuyKXwIHnLD4medIF1Mv9J8iKnVahMM/ewie7nNwzDST
s6MZI/Z2zc5Vr7H59ieO8Es60gO5q2lrdUe/W/rt8nJfbq9t224rmp8c8W8taVKYdMRYqtZvJiCG
0FOmmJLxtROPJ1K0Hz0zUrYKzy55oIF2xCsdoIxQwoURBWl0x1hDtZnc2nmezeuukaBlDT5QQnEV
IiL9yAEkZTGiD+96D9LKQNZHgx5nM3UsAsduiz3lGK9fSKOLCYQnyDl7pNyQqwSVAuK0Efyi7nYC
a9OFRJ9+STlFZoDpLPR2yqWhWDKPfZouZjxPVJlL5Zx71DO2EYvgg4eUkDe71H7snAdQP/Q8/wZ+
y4MMiNcENEaGzcgytE5bUwBU1opcbXd7WPAAvsWhlhzobhAcopLw2mEt7OF+Bt4OZFKggJi2K8KW
ocVwMHqzQcJGI9copIUBvW+YDXTGPFYcI7GnLYCIz32KHOWlmouZusjdveKyQOSNcnC9YobTzKXw
KGqbA+vBQPAhtKzpYsPZ6ItJ7SbL16Dy06/Aey9ABL1P5e6Cn+UgFdvGSgpJ9gQM8v9WOAoiETzO
eu5arLyDYYqWqEZdnpNb82BXgei6rjcI20ZgT7S+fHnTsBo49eMNwVRCFhwh8H2ZJ37/m9Fg65RY
OVZLMfg8Sc3JCGD3JGg6fIJr9Zba+bOn/6UnHpSsYKEwfeQ92kiV295/P1sD3qftGkZbp4vG4Inh
dIaVTiuU8cHz08fcsWTCUZCy2LNm/ekBWimNzfgT7r+DiofBrOn4rsQmu3PkkwGe/A0hxqi8m487
H178kLBYkU02pGIftD6Oyh9bxPpfkA5e/suwls3jLiOXMIvSNf8rsovS/XPBHwLt5YpsYaOBZJzF
uRzbdO487fETLSWCjE66O1m+HUZ0Avz3unllPLZWaDIKIbCk9/pCyQ0ycxJWWv9ZX3ZwIh1f5bqG
pjETwZQF+3BJLrZtgAjFIQIU0Q+P81kGcuQDpGGnLWtH5oUtMre90/i6NAsCeoav4cHAXYDbM+N9
aubsoRmusQwqB8qSTiIQXTCPKhRjmI2jX6BHx0kBAhBDOo+JpPJFqHSy1RAF9NeWPWLQUFnfMDkd
iYm9f5uTS2nrQHeeY2hMilliSfkkKHBhgGLy6jVa2k2sbzAVtBMaLMF967VPf0+yhz6T64sfS29+
k28nh5iME0wYha+Mtp3OwUJjuocm+waHqVAMs2PTLYgWBJP/Mm4B6jW1AgkWIyLwKa1SXqETDUIf
GXsdV2HZwmYkXVT+oBXSJAcnC3+Rw397jQ76oFhOQ7MjE+SWbLqAYX733XQ8na+q71Fwmrd8dXdy
gBnqww0cZ05h4p2dOQIRl3QSePnqSZpP4CgcNe+wnMW4joyGSLBiZf26mmT2NgelA2o1dduxIwqm
UqFIx1XVy5NalPGJn65Q3nAc+ZNQmv+4CYOX8WM7UhSM6untjR47fk0q0v32nFklOI11wwEAG66C
c+a9EMCmmt0y7TnhDOvxni/JYnllgEh6E8on9uSCwHB6HGom4enGBeUgwPBEDEgQhh02S0SmRrdh
Hok+5eVQeh9Q7JsaoeBnV1E1vyNcIg3BMBwPnRp5vsfVsHfUUjw6n1EM65i+PX6lpLfv28tyhG+l
yhcTFH2eWTlmazrgkWXHpfcr1RAbk0OnWH9XuXQ0+kIFJ7qyycV51xaQC8/cnbDre+dMX0JKWpRr
tQYvlgpu/5ThNyBxQqj7zXpy9zglOvBDl7nD+vm1Za4sWRgIG2/aPEV+eFNIwxrXvOdOB6qK1JGl
mSmxyEHrTt6xhuVRBBA0bP9robL1TtIvEINV74z/fR6QAGEPRsKStkECT7V1bMu+cz4zM0sjw2Uw
FP+8LBmULsN5rKYhCpqBDuzn2/Jkg6owavCyNevRwADLIwASWz1stYdpjA4kpOeuzTQNFkUl+Kgz
UOEzBKnkApOduSbwbja+2u87qpiIr1y4Vhec+9zMyM4kFaXfE6Y3uZrM/qENn0WAf3ORNjMlRZY9
m97FqtG/Id5ir/BrDaz+SYL57dRqFAp9uB1EhpjyZwbTUIh+sK7rODPduV46gfv3aT7/1gdsoBlA
RVHpZfflghsaF0rc1b8ICGa0OoDJ/O5OyEvxBm5R+21gaqMgjqdyBCUYDJ+OYftFVUo8cw7hw9Zq
BUOFuUmHSXOtec4kCO8JyIM7IA2VRogfeBAncKzhSQ94BbU05s1ey2FtiNC+4cnyV7oUisB6n8EQ
dyfTC7jNvS3fR26Lfsy7Icf4LALIqHkz25NUJZKhuuOlzY7xprRcKfau6SLrQne8RQ/1SuDwDLA3
XvO21UUGeAZQoUhnvYOKiKjk0dHUzTH2s4dNQEMGEB/d5DvAbukHIrSaC0dVpgqnxW2eJ9Uj147e
ALhR0UM08FGLk/l0VL3xX6COpElMG2VuAgHdOgCgEd4c3oM/N7U2ybcoPPeB5Rf/XFrvbwxnJfU8
wI/s3A+/nXy02GAT8agFXEEgEmZzT5Yh2elb3AJ3tDHrWgRkYWj6+LHLbyoBMn3LznIkwrrb/gQL
vfsYrqQocp9AygD16RG271vuugK3ui4vOZokKfKsBz85JkI7dQLh2rjmcztQa+Oy+J3/+NkZMkuU
p9JYepQsOHdW0Vi9DsIuyuomSsSwsSTLe1rekPJzMpmY6BF/ep7/NdagzvEZ7v3xm4EiVkHxEqMa
SA/JPRl2vDldxvqZ18nRlPjnL4A3FIGSIZcntAslwmEt6eIybS4jDUxF08bqTYKUVq35kqWiW7fj
Bza5UWZkC674tHwRQGQqK/MDJWRs3Zk1Z2RrKZl3ThAE+RqjvCjWgHRwY7ER6Sjfoya51Ryf1evz
jh4a3QtnW1nHMcrE2Euv3xcZH2tHnT30FTLAt6RycR6Dtr31Qzel7MbE7zMcOiWn9OlfPM+hSNDx
B5498thZKz9HQlEAxge3lPUr7+McL9e/uLjnPHrwpTBH2PclIEn28Pjib9KWg0HMHLaGqIa5iOJS
L8Pxb/A5GVRUhUE1F7XpyogOS2e1sYwh4WQ5S5CriMO82ZSQA1squ8lcMyzFS+eezHWSqWLMeReI
hFdhCiI8Fu3HKk2PEgRKtaVxA2iJdr1iV938iF40GFGiC4V5gG909iXBMHMm1xkxCLXFKAZ1LFfn
c/QgaCRSfxX9nEw6sGdpsKVHiXj6WfD2hUzTo4191rpVCyktcs+4mECq9o2CcHdejkAy8xRjYDB5
yAWCDwtU+pxvdT0p7PKMi/rnGBDqKTu8pSfM9dCE6QyFl08V0s14cD5ziJKah0V3XfU+R8r3D/9q
0r6GhN/m+fKsrCL/pNgpsF7eFsRozqreyhqA78d8Pl8Mkmdxre4OayHGsCNQSNL9wX8DzhjuWDah
eRIljzouXiq6XFZUX7ToWHLKVQOEjFP83DfNVIrEnvFTGQL36ARtPfSd2p8DEG1lWjDUrZnyyq41
l8IvoJMwocLElC7EahBTZWeAISsTxjYqxWJAFYrHZA2vcBM97dJ49dX84yaaSkqYzKaCUHBK8nGk
b5knKlvp97CnsC+eCFhWggZe5pcYhjX2Yh6IBM1IYaXPYufI/qeKIGGAY/tc+Y5gqyURIN1YUYcH
Q7pzBtUCAKpdW+sMvFqSk6EDt7/NidsU075UcPLa1yyR1Bhpwoo93pmFUzkehcweV+iLdNvAf+6K
SkhFrDGMPFlLEWnMt9Uoqa88J2RVwIkK0/R4QnPiL9id2EqJ2M9wtpfZwVfO2dPswgtR9t+00cdJ
wyKG4OsK6o2Ao1qSxyB5dc1lzgyumszOUvzJRzMFtMhorIx4Z1L4GE7QdrThk1HodcS+MLAflMkP
tgHLJEV/ZpfaQgr4tulGgFYevvnhRY0EAhp76/75/X7JeJ9ifMyYJmV+G0gytF005vTOzVLe1RwJ
SoOwCdBayryJKBJmSe4gqz0U+xzA0JEZd43/Yjd0aXGwkhbnItVZesGteTz/JeDeV6bEetdDiOp+
19hrDayNHjcyvGcPyMjtvz2o/7mA22BxGzUObBGyewg1seaACJBi7vWST74HHC1z7zro90Mn5/xD
yaa7OlsdpVpSkK4ohJAv5NwbYXrYtLdbvgCToOtuRc2Z5iDxvc8C/Y67VRo2f+q1U89pYaafMXeC
Ktwa5ozZrG7w3WI7/HsmsrK4mb/EAehZdTCgfdVWBPxdNcqSJBxumb5NHRgU11rY/tqZjBPbr6Ij
qDf52ojM/bMdMWXtXCE7FeYDpCl3fL+ZtqqQVAc6SubBcWENhC0MvCGQHZhBdZMKSzl1GzlO0XTV
p8zMWccYlfBkZ1vTTTpRitRLsylqHuPj1Iu7BDv+gO7gHxWVgDeP753hU4kKWAkETQdkeXBV9s9d
QFTX6LgTGcFPeG/hyexvBcpWYNuRqnXYCUHNhOE6GwgqbKf5lKGs2JtQunNbIKCgiYC9mjZWTuyi
d6JPwzOAN6Ua/H84lpWl7ViZ0ICCCeb6MRaWlCEOYi0FFJFhMRo1IXI5oU38+oDLVVtUEEzQ/f40
M8anTCM6DhgMzvOkYO6B4iLW9OX9xS5OKu6EEW594U90vk5z7Io82NVX4fxkRUD7J9J30v8c1fZO
iK5lP6KooQwtTZ6Q5iEm3Y4YUIwLXLDTfpOSnra+kiopdYHa/JH++wWTNygs485lRnJW2tGWkDYc
zdoDH7OGmfiVLGPmhM9iJoaYedzor0YHkKvOsjN9mmPb/7PaNFti/B3O1qcxTCP0IDlBxgBclcR9
GSbwyITRtK+qKuB3nbqqjhnbG0afvhciPqDT9yK6sMZZQGH3JQZfMD+EerYJIp7CiYZ4ujbAOUWG
mq/wXeVWFQbMMQaFSyM/2hK1dk0GxDIo9VQrWqWhJ44ORP2OrdIZhwnXWQuxPZmM8FNd9APA8MQP
ua27ehx7VHmktf/vOdX/mzyBP9UyRvCMcl9n9GZj7qa5YZZtbF7LxPHVvPh5ubaxd4CWuidzOgsP
pdSn0Clw0GAC9Qy5fAgSm1HaX6coXCa/ynq0IGYN4VVVRaeMpT8zIUeuVZiEEDkkY5D5ilIMfSSw
ssd8HBk0kEKsE5nrMnrgm/01yKOu0lm6QB5MC5zA4ejmF5LG1XBmxfxxnJ3cjBK0snX+WKnHkNMc
g+0wJSwkvXdqLf6ji2b8isoMAvx6VA6eDZINSTocDmT6qWFsVWI9/dsPggVXL7g+Rhk6YfpB6yjw
w/morubf6PV3pMAgNABoMiC6W+F2ugP4DQ4V2VxMrqiwdRqSHD5WgUrXeoiSzvdSvdHpm1LBp74g
m3hEzO1J7fc5tXUZEJ1FNXsY3JqnwAkqvBOPQHEr78p6JrIssF8xfrXdEbpqiOE+0fxnODFo0bny
LN/P+TZBYXyuFV9iFgxFUMF6JLbTq9IR7onz+8ngz5IqpKn+1o96qE01DP5WCrQXZ93BekNPEq0g
wZumKxFq5TNxpt9XgbavLeD4S90P3sE0SJK/8u1iRfoMbQ3BU7xlHbGQQDoZNTAfnMIXSwRAQCEY
iBFmHk3d8xRiDFgHGdZmUTyKRolckCG7UHG9SAMS7gYTRQ4RM31jSXPURMugpO7fyUp947o8InXI
iR3GaxMsDzXWVdchRPurxhm9P23jZ2LUIE+Fe8PDuR8VSwbZohPRmm5AonY+MqeNloFutYUuj/LH
RbUaoxR3HkS46JT+uvJZ38sVqLzzoil9uOiYdNIEL0H78kvU53sFACmXyCw65+d/pMx2Vim6gYz9
sEidzZMW+Cfgsye2aWk9u3pszGLBRsi6WzaZldDlNQxIhWvi8s8EDa5O+MQM+GFCpynN8HVxoL8J
bllS0hTSxPZW34pNBPgLV2UE4dEAFNECo7+BHaSGb/LSaoTenx2SIoX0k2foj1LgaLuRfICTnP6Y
Dwgzd+RDzpgbNywqqFo6SOgshwk6snVN4nb2BortKWlRXx0KvnynFx466mIt6QHRMccLDauQuzg2
8GbFoiSvm3pmBwkMM+Pg6D+SynUrsKIDaxurxFZtpgzZOk9lX8DvZfydilvUqGOuA9VcitDeuj9l
BA+buWGJdzRVr9Vgl88mifHiuFLJKMUiCAk7LU3TZ3jNsrluZzbelD7o1+kEWqrbveSPVajyfBQS
3L0SuAix+pHNELJRcxaZ43RqxTrsVWNgwLAW6QdTZi9psu6LdBXJVZHhUBBCRTl+wv7DUvTIyWGL
es1r1gUbBRCXMlzNwSrvU0sNrEAJ0buPHlMyks3jNt2y4/vXoSowaoM6BJlUM/GRqRSbe0tFywm8
qZNyTpDGEYBQh78wauUXo+tcxcrmy5uANPlYeM+neRk0BV2KIaOn+5F52AhNla/FEJhhXvkmh9S+
IVvWatvtQSJVr+KPeeqxa7CQ+9OyGoy5jFSx+Y9la0Je/bSw0xIz3PLq7KQICx/N236lbYZIyfP7
e0qzgRUt8u2qDw9yka9p9ZeUlQkh9X5px/cLQZRKOlkK1jTeA5QGZksrEyJSBcTA0nrBWADIbCiE
c/3877UYc6Bk3zkq6jvDKVsWmmxatSBLSblYpTsIDHkxGT7ebiv6LfYwVZ7A10jvzUp0HlAKssK+
rsDUBaNIvO7ehAnjBk1qByT3WdH0RjNn7pBSgHjru2TS07d97vvycUNpEGDXIoNv135s7IYF56Vn
pRL4F3tQmBbEu1okK0IurqE9PAymijBCdkzcAYhqNwnEKd15HZd1+Khm6UariZ+dnkKO92drg9tV
mZMxTnJ243VsDGWXznGl/6dMKCprwB4jhVN1hfQB7yK+WJkl7fEHYlaDvUgqhccPkWhjl+tX6mS8
SI/y5zztUF5AKNktBbt/TktWtZseX06GnjsRX/IFlzsUab25IpUNUTFEvmUvrJ/Vweu+Mr4YQ25H
VENMJZ3nAJ2/jk+4+loFgQ2/VhKz2k/t8vH9QjcB/YV0E7RhkpXs3nUmu7/ieVa6XG4yrqCMRRBd
6QaaP4HslgjebblMFLdahvSQAcPfvXQsZx/OpLjFds5s5RKnKoHMAXF5INNM2EMkIiFi85L+VH8K
atpgOzzHiyrQVW62RKaQujLf4BarN2n4oTugNLbECtARXq6wu4ptpCbXXuSiqGDK7DhBR7vBOecZ
DqF3kyu3V+TZkHdfM1n2l6+3gsE9nOKa8LTY+FkmSopxTiv214lJ9vZtRjKj0yF4WDSTuLdlUQR8
eApH8dVjxFEEXEI7gSSzoEQbOTcLFuAyniXix/P6CIRJCI8GAx86DzyTI5HZC+DNiNyA3Mykvzjl
KBKEjgp5jG7Ri1nfC4x5qtyzytJACjm8Wh0c77wRhA7qNEN6sOcpZcJrcsIZwR/lodElXr1DFrha
Q63bi0zZrET6IWC7Tw9etZaM8WZATMqphaG7W//+iV4BIgvHjFNgnS3+OnZazIC3EQYRDXVWmvGL
uqTN9YHI3hr5jeZiQZFN3OaesR5DqscYfDzK5e25h1Z+cgb/banoHAhmaQcehFBxD9VQQbUGHBsF
8/gZYOCuHpbU4otUxJGwpTPbvfhpHcibntC1TpoH/oZdlx+Jj6EJm9JjZ6JSAT0Dkcl7K0nmtcmo
tPxQ1c1btiUt3gdjwsJyz/VMHvfF1XgCtiMV1UfEivaiwp0hPWmzaRBdMYeWIZA4Ty5LnHrecFiB
lASBlCo3p8JQ1Ujv2aCLuYuwegly45VBjULRYyn8Hayj2+ydZl6TBgCMggSmtW3gZN+VFx9sSODF
PwzIOIeEmkteSj/0sRYJQjrEVJr3iCXKm2k772f7GcoDq4FszhJFalfv+um81M97kINC6UJgYrtD
bPkAbteg5Tv8mgZH8f5uwEhPRTVdcOJfeER7Z4XhS1s7juh/+73lLXg5DTYRG7CLFI5RsB7Igy5U
w4psMlS3USCw3gTfkHksbC6m/Fun+4wiMxijF8P2B2dpAqpv194nMnrmLuqaCUZqPfTOw9jfpIQe
qIzlBH7QXwZOMpkG9kcK5dKwhPSvC56jsVqlFXJn4IXAPXM2Tznrx6pJZt59Fxmr7FXorLuVyjHB
u+tRDCsdRR+wtXBHD4f4GbRQp4v32V0VoljxyV9YznjTFXonRE77+AXrf23TwzWcS25+4GVZm34/
bu2ea9+ZChdJDxpzyxNCTA9pgPLVLix44prJNfOAapVzJS/MU+b37mLP7puAnRyCtcTr1A2vQSl2
BzIZXipF5dT+dIXkBBe7zoRBWErXSKCrISbrmVfNfWmbDOrTe6AjMatocxgTT3kcelqbwkZGf8HI
F2LZxtqZ4Ca8R+punEpjaCnCBieGywnUhEKjvMqbTazYoQa4MkIEMCovTV1EdXMZt5fZ2WT+B/P2
jOK83PQZKDuhaKC0aX5BJMdPdzrzBgOErVdTOO4TmR6W7DzVHB/rkeIyN+F9o7yyHHRztflyZC7a
/LwdBFiTxL+22PGJhXrtHjEVtIHrxVgVw96NDsRnD/SzRDHW2/3Qr7VI0LQVGodUGfH95Qbuw/Up
F3IDfz8wuIWBTIDZcGfNK1ge0ITnoStX9cvyCFRO5UnqeNzoPWWfANJOaodtLsxBh6mcOiYOtS96
RWFl/AHUk7HpRImGz7aJqNqInHknT7hHCv9ne2ffqOkr7DCG0FtBmPlGmYsIDjShFpB/aB0s9aPf
RHhb6HPvLyjxPCncPpbvEwhM/eJETT9MNN8LdjVhvzAT9OIBls5A0ugqaOI+Eng0tmcV2Ddx+4w8
r+fR7VQvdpcNE5UELuqZs+LOoNJzkAJNLQxXWiecC57YR9VV/Kr3QWNL4D/gkS3CEud8f+Rq6ZIa
FzXidSGStpDyAiqNlQB2BTQOV4R+IEIdL843A9fIDAQmzw31omtwn7ocTbDf61uFrtBw2xDn1IT0
cWxtfZ3RDvIMYwJ3/QH3dCHw8rCZFQ0nvoJ1quSocurjo8sfrdRjeBMKE6gxocgQP2i7s840rXXi
2ZqD3ga9MLO10EHssGJF8yQIvg95DdcBMl32LQb8VbLCoQJr2ZoERZSPsvPh1TTg16TWT8nB26xD
NcQByh2yjOSWw1ltaNVHGO6CVFH+QAO2JLP12m0S7/xNkqtLPEt18nKqLdsld7PvCkhoXpPEIPkq
wR1w3HpaanNhXNwtJueCITnO+GGdoL1hxhKSmu44/6ptKPmTS8QPNKcCK5rv/TaBAzOkQni4wJfe
bGNZVFXfZbh3206DwVKIgLtn8XNZ01k/eWHQIEXtgt1ecwanwBEmAPTwrEb6pocRBm5iIGligGIf
Wz2uLw6mQRc8caMACxew9xISQwGVOkH9KoGUvnmf5Ym9b9dFH5fgAdK+LEvySRlN7Y+VVXYHShGQ
KT/fF/5QVvTb+rI+6LW9Q6UR3sbDz9fGkYm7822H7biAuQYxX5HX14Cu/bFNtXBT1Kiqd9F721g5
UZaHBYwG65LDTwiahSUpTWw1UWSHFew+K2Td1ILo4DziBGYRrxsg8gC9B+6y3UR7EnHeFIvGSrR/
q8znJZAxSfNqdaQsYlOJiawGHhSFpWBdsUJampYSJOzNIHec5TWeKmYmHtsklM0+uPYSCIf30uKk
t/X3BnKQjIqKt6lrTATl80PzjLfWDnyEnlSWkU+DayrdGltzrXklzS84dqMleWSOj0+bFu+MgpBh
wnkMo+0T5YmzvWIskKLsv7NbsXYPIpch+9zPSExHELuuMwBdTJFt4TwG1qr/f+rzfPeGLKgFeMs6
VUC+LosnrLeCNYsAyrT48J8JG05TXYfLd5UR3SrnuAWa8NG3nH5TqWApkQ7QxHU2gF7NAr9B+jTa
qU6fGzpKBOq5atmzQ8lvE/vuwBvMNyD20L5ehJNe3rONpeNDrosuqJcYaNnUNr4Zu/kzVBv1A4Dy
bYPxrtAwhoHFNT0U4W1l/9adMTTErWJh4rsC1aCSoed1l50Esyr40BSavC+GJ3tLF3miJXvyu+Qh
Z3pm13KKue0mJwwhO3tnqrLwFC7/NexIXboLj+J2IQNfpObh3jxKlp+pnlO09YsRMQoeTcTa1Ahd
cwwt6Z6qjs3XZ9FKCIJxniZXqFRaNwQs6+8NKkeK17QPDQ6kd6liOSaCDFd1/XIS5TlO4/xPn4AS
mTXlksRoWMwPuanGX57ZliwnAUXoemT9qqWt3wJC3ha5cGsX0C4JjNpTdlQyOiP/us2+DzKerSiw
+NLr/quwzThazLaxJZZOVhOAvabJA4C+67rnAW9KSKZrJabeHWVTRyH07RASGb5Ky19gelsV79Ng
MnEs3hmhXK4M2qYpt71IHheMDEHq1c0yb0rZHhoPfgjlyqX0o3JqASjgvcDK+8evUFfwhNBy/TBu
ebWm/O/SzBxS9r1kdeuz8kqh45B7bAl/if66nuEFfH/9FsgfKTMeg0GOj7mEg9wteJloX6TFelv0
sgG2Cgd4i3wMg3mj1C5daVrb2gSGjGUNi0u3Wc0GmkEZ6+IEhv2rEHUAu+ELb6noIm+kD86An8nB
d5ryC0vy4eDC5l1fVtKOdqHPQtuWKqMwJTGUh/t8t/juuqIQQTiRy8VHU4wxhpwNrnJ55Uf87DEu
YuWeC4YL1L2AA7xlpq81axNon0EbbRilQKy3fB8ZuF6L2mixCvPbcouj3ZRDBs1ul6R+XPbSBkhY
DewtS2S2Fb7lmjsFJIuvEqWke8R08Ens2rf7TDcYZFqI+NH+CTm72S1Tubl+iZE4gQ2kNP7lMT3W
zfMZIJrVAiglQdilrpf4xlFXUxqPWBvmgDH8UVvXfoIUZodW+ulieV1X9JNen/3WfpJ3HwNX33PG
rOAkG8NLheLMzAYMyk4rSefM0bpj3Ql+0BqSxdOYWOzrnGIEW5ZljmDQAS5aXK7L0dG249XwA7As
tL5cLkrzv8iz4OezL3Mw/HDmLmKvRtOCe7y8h1HJjm/qVQqQzEodscIPjZRhy5icP8mMCcQC8Dm7
5YuNYKmy8M00Gl+nb2A8qmRb+lbbk/iXW7X3gVNDbWNekupanFOGouwYq9ypprzAKPh1bbDWc3rX
7tqjEymOFH3C5/v/UjhUirWKPgpM2xAOdhW1dJJQt3x6cj1Alu++mfq2ZcsfqhrliGWTr6yvSrQ3
kHppX6rnLHYBOOoXYIs9WpLLSNj3QrpphopN4PNxCFL0fDTEzJuOE91vTNK3ONmUZeDxU4Xx6LI3
0sVm1DjxjlMKhdOCTiO/AVbcPfSItPXc/CgLdZTBy5K9+u95t2gX3sXyyl8qC3YLqbrttaKXfJ29
4PA9AaB4aF7OvIlV4OUzfbfNksu2EZMZ7Lad7Ml0ifbCIm5foS0fQ1NjlhbLHJT2RVTeFwTpXZPe
mW1xAzkFHDHPg66VdhF7E1KMRhQZIRbJRmqop2p5dF5dUCS3JEjLLNiD7MId+CK2qZckP6SlSLV9
QyhNMQUU5We1TMwZOvPbWQCjVrBx50m+dQ1RU1wv4tLA/2gQH9CxYXLaD/Nfs941vmja7rXC7+RA
CWrldCdB8DVm9x2Pyw3gTo/IFlnkY97Ryl8WEPUToKSXt7ORIdgAWFahlTZOUmhIev9lHdHYbY9t
b0ybd0tmYXx7b7L1BAv/cfU/Li9DqVtryPprmiGBzEVFAtMYEXYOD6CRArXwJeZtZFwV0QerHeH5
VjJGN5IDaT/kM1pVD10+C4AHIqy0yvwJDohQ0Y2Fh9ncieJTklrUBMVkfNqrcxG8FslMEYzMDvE9
pEcu0M8vsN1MFvBHwo7ddUDLaF/bzpOddKgpnUrZdMtnt+r/5K49mytGe4xS3gU3wzANQXq23zUO
ptLLhydEOEswtfo3jMIDrZ6NgpODOftz0uFSAHE+aSIYJ+9j2NbmC1MPcHozVB3nO3cYz2/JMucT
QqoRV1ASD4bflDT1amtq1VYYWtojaQ5dHwZIgQNt/w54IOVN1Eldj/EPwuydiSZ5AKquYGyaNnBU
fZyrSwd8x9U6OczOxJouwHfE9nRuZt3jtguvgNHz50QuFIulP6lM20ZuTwn4f3233gr2g32eX7i1
PktLkYHoYTS6TItPAOpkG6nuH5d5yHzWuzLYlqDaVO7qV61TZ7CVEHyE1iSTdlCWMWfjulqw2WCz
qQI1ZIjSq3LIUBJMTzNK5Pd9X2Z9mCTHaVeJJum8HwmH5Q1jC49dONZjXnPlYQQF6ZVaTqE3T1UX
OMmAYsp0qYF5Scp/Uoee6Yg5QOJq6uTVM/QEhjF6rPAxjW0yhcBPHymdCvU2UrKnvKM4CcnTyzYe
FbtED+/Hpwn9DGV9lXm3HXYhCMU57QPPD18yMuymEf0Wq/yUgO9XMYJtznY9QYZdyh5ZLazjA1ak
EOQ11wzBlTPZGaLmnAFuhfPCpNVEzpzGgjkhmHxfMfRzWormnweUBQT1Em/oO6pcv4LF0W9sizDy
U43DXLt7nZpN46YJvZ3suFDGsLcjRAylE7tWJEpIbFvzEx2l5oYm6NQLbzV960nqniZw9VCwWud4
+K+lAdABmGEF7Bf4a6P0PThKZMFwXxnf2cES7U/ZCI4C2KRs3vvMLpbUaXoRl5loMi5oHW5rcJVX
ShDI5Hx+tWvdsw3mijKe93Ol9lD/j2mjtO5C6V2O7I/0+aiozVVyV9Q+KvnuFuyNXM9m8Vb+BmXx
C965DiCRk1kg4PoVHpqe+9S43BkT/4SeBDuqbE3wnXh0oDnTjW//IlVMK266PgWEa/rjpWGKrtOD
dYbM4xdVjUvDtWzbRXaWSmedc8iM4LsV56D4BbSqTrv22LKKixECK4SKGGFEczQk/PzEZIXvnBdz
emGik+VE0EvQSj6x8so/fJC4SF/HHdJy0mUD0mF0WaFD6oxzqZT34rkxYd+TwAu5d1kko5ZeTPUQ
w2i5erK3oxyTGl8dcHAnPbyHnVi0/ILA/2NeUlkCdt6b8uPxPFy1w9uD3i5dle3A+zsrPPhiOj4m
b9ebY78FQeG1pplqZtwMycfzKk/pxth4mxTslUNBwHqrg9ybSyha58ODU4Z+Obtr2Eb9wGHFbgnC
DiVXPVTfq/jyIBJeWRNzmtyXUsaMe1lXRvJXyYy2pXK/a/E/jqvrPvcDmDI+6iyaKCJhPHOIRgyf
UE9s1NtI9CXWR29wvuDPWgcUnLc6dJr2jimgIzExsx44pjzozsXQ4Pq5jhasLW7zY5sFOkitu9ZK
WxSJOaG0KoDuOdXAQuOmeNyKNN5FFTfTz/jKyXUIXIQ8j3TIq7EsDlEEqkUmyowb45fG1qVjiS7T
oEPSx2zLscmvPS9LFZEKBxXvkXl7NF+BMODNEwN/t46XcWp+GgGzdcq8UrxjzUIElA6OooKC8+YS
FFD9cIU9UkEf0/RTLffnkxoZ5CitB5pYbqtWSJal8/Jfj14r0OWynZDZM/cRKRjns2Lb52YChOEY
e7qO0BjCMq1agDoYmp5aDOvlPFjQw8BLeqmOaB8zbZHrMNWZtLbhf73A6X+SQNnkm0aN3CoYuN3z
uYgMW9Io0dioQngWujlKKfF5IIc926pyVXRu4JnAFLmtcFFDT1huMr9Gbf+xocGAJfGbi7IRcuIh
nfIxUU1qnL8CQjUcncrI5Veu7cjUpHMv1OgftwXc3VUqrIYaLoSLCn7O5KeoR6irIADjpz/OdNMQ
3rta/MBD/GJ+eTbt//IROruXLNDbcuFA9myDtWsZsAfmfBfsWKIrpkgNpnxKKi50vu+Ixq4a026j
cOkTXU5ucZ0JytrUBPMNh5tUB47XVAEtvd++YzbWRrnKeNEB2GxlGzP1FhNsy9nGSDG4NjHSidGh
6HQ23qpH/SmCUw2vCO9AeMJYEtNy4rc1xshzUNDeI0gEz40SMIFceGvLxip+ZPmBl2GaG7fzG8W7
2/l75AV9E2u3qA09PejkeDs+JcEdeLOmmqwLG+2zGrSm/9IS0dmQmQWu0KhZNHxkyqwKulbgtz9C
ihv3JvJa1tDWwOM2FcUcd/q4GrI4UM8FUK5E0vKF0lV5h/mbpMHT4yPkRvYN9SHHtdizDPCtZ5Fz
Z73H4wYiz0tqLwAxIdL5jP9QI5VDLIkUJZj7rAN6t5ZB5LfM9LhiFcg//KRio/Lwkk4zzlMCw/au
5U+tiBKbjkLGjyv7ADPpGzBGpwEgi8n33R7zQF2sgHzDMwlVubomJqlTh+DCU71xqwjdG4R3d5LN
OChyXXzMoQrzAOLVP/ULCxgvwLNRfI77Bx8sI7/chx0fMD8Ccki94CUoejT/Y0mx90YRWr7ot7fZ
6zJ1WAd76mLI1uV8sXu8WvNUzTxim+iw84LfDALLevuUKT0a1568sFgvq0KUzGvdxw8ZzmLApkIm
IFmpBbLDkG2hm1X3+Zbs/xVN51U9AN48UwrUP7TNpXY8h2cuJ6l/Uhw620HrxfmOjuFl97Vb1PPl
/DBMBp02BoZrptFlPC5ijqU/4DprPlMKWIrl90RGqPXhMhCJ0GWKcVjztTuacMBCR8U0zPVdVI0q
ePrO7NGLr2GmIsAKlhu9aauoE5dqOXZDXMmz6gvauHps9oMuC2PsHjygZBMbU+GcIf83rcP1FTKI
IhJvEFvfwdeul+9lkZUu37dgOAe8T018km76zvUViXPHRUwRMD5DRxv2YwHKNT/zw0t/ka8QeHw5
aIKtf6JrvI83lhBTdEhp7K/QvYGjSzr67+Z02QFpr00u3k0TSfvdz+Djf6hksOsDSlC4j/FHoovQ
kalh3aKS+8iopl5vYmJFLw6/l/D+p+TQSxTW2YoLQa4goEaI9AM59PVjMsLFYty7G7199ZVN6K4i
LocJZMDcdAeDl3CSfoZilCsee6N0A68f6IzPMeMQbduLF/fScBlkkEiAAPf/WGUTGsW90xXwwN+r
PcB8pSc3Ph/KjfcOH3WC5knVvCaVv9q6DGVwsCMckmtFZMAIL2UEN48LXtVApNZmiLB8vt17mDYP
QEmZzTjeT4OIyWkA/CoII+kppCAqExa/1Q2ZdibBsFoQO9a2S4HYhoPyDAXOUacjqkuHKMJ6rxGw
oWRJSXl1pKluVpB1OnBFLVRmhsqjSU+OEIg0UZafaDLy/0c9xD0G9pxNw7k6RcpTEK4HfjHFzqdz
b/kvpC5pCvg3iMysqd1xMdl1OPRVb4HxmReZJMo5gPf0hsi/b85sXoOdG5/0ukru9o91WzsBGQB5
g2fUpPOLUMLnjV3sCj0Fe/0/H9e8OydX/We8pmJ94b2YJW/Ai1stySACrv3wWnp7V2QrMp0s3QWi
3pBip9na+OKoy85wbHV3sbi0AKFSX5ZXfEj5H7pJV97PwNDndiHtvK8cih5TdVSgdThwMKPlHu5F
YruvURXyUwHK1MRQKK/+SFq7KVkqrmiU3ce7dn8pCG0n+xLVrWg2bVMml2mRUQ6RNzHPeO/KHc/u
JqXjRS61fkJ84e+OuagUUNGRgp0bnYc7x676THvhnh34cqtPaxTCL1r1jTBQ7ZuCDmKUYRO/OAFp
IbceIii2rrrzjYCtoPSjvEQmlyJkyuFsq1mpWOoBzL2tQvS3jIn/4xVstjz3pTXau16CM9hnWwLE
424ms6nZZ8QWqmsf4lzvOPhOyQcL2HJ/U+oAU1A2ZpATq1vlKITohUarY/hV9UDd9y9QuXWfiaXn
u5qfC8PCy9SriOMOweDz+QVoGqZ2xl6f5OiUUhfNGjYJFzrN6sJpWYyG9IjWFMUtehdFhOJJiU56
ssU89SbivGxnlNe5myn0VIdW5k4gbLHFEgT80TG6lfT5NxBvxh+MNo6p8ycoCBt9T5GafBlqdPNC
IfJsOV6zgehSfVo1pi2w80JRUwjn/AgsE9XQYEklCvLzQ7DhQ1nRsy5F9yUggJ3NVBMomrfGqkf/
ARF2esAZ706OoEFcId9LvOQCT0K+ZDKRlFL4dspzCTp5gbAD0CkY/2JzxwdzXxsDDd5VzYZBaTJC
OIlfzD5KfZ00Lof07sBh6QnjeodCUXP7hp/+IBT2Z2m8E5rcDPzT+7hZ+Ye3eQYR6jzsqrEoH1vR
r3OlsvR6SpUQJZ811CBthk8Ohe1lUkA0cHEb6nhg5yhuTbbW2G59ILpO+5bJqa6SgE53anDJAbC+
dX0bUAken7hJQ5f1gYGuNCaPMEprTTBzwjPRvrTzmsPNIRL9rQHHsAwHvFUpU7EYghKSgAgqIcYM
bUyjoiJ+78J7GH9iFgHbolGrl6HsLn8UyEFHDvQdariCW95RuqQfzxEtIXRt/vv0sG3qVIOp//QV
AaD6Qh1564ZyMS7w7O6WNui5MO7pJrOmmk1OD9MP5haF8NxY3lD4CFgHraEbMrRMz/0GDmxVEWSi
QSL+k5sWIgxVxtz/UdAMTCFOtvrrTgwq0IehkLcbexpyGKh/95giSMwhN32qgBxe+9JEzYsH/gLL
loJSMBXQDMmcQJ5/iwwDvpoRJaB5g37aCtwlBA2ud3+xbgXlqRx4OKxGsjsjYK6sQb4JYBcAIuCA
SvxASMlN4hwzIrjrGadqzOwrMzwcywT4gKTnGrGaNlyE8gf19QvcZffikehtcUF7h1Yq9rbpFa3c
QYw95I9m90OelL+UNp0JqufpcJXUbEJyynYWZiqrOKS01n68eipgGJyLdW7srIz4PgoOfm8p3wLY
z/Dry4ACGHVY5EuBhB6aVM1Fpn44p7HCZBqkEGFzbCaELWcUTI8inUs6W4aClHjQDdEbuwEpCiXe
sDK4tM5NMMLDf6Dq6MsOkU2Rhuk1AbKI2Gb2xyiIn55PEWCZA45U3Iqb03/1YiTCzGS1Hdaueqsy
/HIasfc46G1mFALTdM2VfjexVaftRWyJMH73Xp7O4xfJPKh4v+VxlXZBSdqI6SrEhBBnmNsHtPyU
2fVL7gY+mvy5FWJhYATATIOj57UgeWaXr/5Vivb2/2O3hVPjBzzsI9G0gXVlB3cgO01+wBlNT7Kq
In8Bhnq+Kw13gwAatQVONwU4E4g2dF1u3jIyXTKwchUG2QNHac4hQfzJ0XCt46o30pOcko6GYn8w
26hr3LA1RkYfUUrzOrQb5Ia/eztyxrNGyIO1++rSjU7o5+AsbBy0VxB3E1a6Opf2pGOm/gT09Kz6
NS7LXUsUgz6WS+Njl4/4CRMveHB/TlOZmTo+ovf3B+IB5DVpEvcKIxk23Z/pBTDkZSRpgA9MBcej
dGWxFzqkNwEVsar9KN7BU30RpQ2j5gISrtyv1B6iAI/bOMGATXzw+vRX7KNQEtzqx9Zf70Fs2WpS
or1Pv3py8GxazQK9sahsi7t7EjQVgO6M66O80iOz65TzYU0/7hnAPihfWiyXAk12IUF639uYN8T/
xksD5yUht30T4CmuEkr/SY0G+AVy3LFwIVzBy3sr45FWT4sfbU9mT3sfZrCv13Y0AEG9v4blCvZS
izurq/wyRjGWUho427Pam+pGPGBez6ilimuMgrx4a9XLFxbJwf1Ok9CBqOsdeVne/ph66mgK7R+O
pTMN09V9E0y9jpZFfpSXx7eBNk8zyib9igy8t/xlRoHGlBZdZ8zg13KGkoYti5mpQ/VPk0nJQzwj
Wg1msqla3a0tUFwOJMaigqU6vxQbCllGIuYYn808o77ludz/OXYK/YF/7aYYWPuNr31qESDfrLwj
Ty8zXOXr+YcBovD94WXU7sndNx3UtSx42RhpYcc+9SBrfVoMM/DWx0FKn+gmZ4sQ7jmGfDMMViO5
nFODRD2wISjH7femtBTcW9iN08XYixgOt9ZAVqEWK8U0/hjR21NPk+e3i/bbQlLo33cikKdF9bxf
KgFVgW206UlQA9rDa8E23DanrnqyPYhIN3sH9W0OWD6eut0HcosoBW1lhY/TUQTF8Llu8Oo2jq/1
2mE2DhDwNEY7uopTrZqrPH/oDf5u1oDbK/yOsIrexkQPxZUKC5HWkKlPcTgfJj3BQAb3NdFvKylJ
44qze4WO2QsawvBYy5dk1jpVuKbETcFn7FmPCZjaY79Sf6++Dg9kfgirWUjhjsISfjKTy5uERRxs
5Wigim1ugS05xSAzqgOPFaWCinwTl3yMTbIS0XZQbBBQPz/ZtyPtBecnjdsrAljpWjLdUCuhTMjv
vxO/kTCgw5Cc34NfbahGMiWcTHnwG6cM/7wNtyQ7aCocXTtIOKB/VMLbMe3JVriDbhinqdjptEGh
aF0iFjbSxOvYtJSaHOsq9k/oDa7nC96+7gSBoymcW8NIAK9zYqma/93SChkEvFvJj6nMsP9f0GSr
jvXdnM30/dH9TR3qr3rIimHAehmInAP2mXSFsmm/ukMTC27D17QFXR2Uk7qHlTA0XasxSq8Q8xt7
QP9VKYolQ21/ayjEtv0bg0T5AjqOjNbwKU9s2IwryFq8IyQ/VWRIF5bVKixeWi6MuuF7uKKGQ53A
A8noDTfZF8gCRyt+HRHI/aPV0eKflVGYOJ/yNCmTg3kRdllX9mk+k97Pgs5zCifJpjgDk5PXMkZt
CcRTqSFRkNQJhuXGj22RIbO2zAkeMtNUGPS0uZJT/eDXKTr3SFI0x0R7G/1qtW5NOTyyUWHBG/k+
NvVPVXIWMNNCx1iVJPzeSzAC8SrISvY9s4tapMr7YDsOCNkGEDYJxroxdc17TblTuSE7uYqdNi7c
jXUo1BZwmT/hVcW8tOjYvsrykVFL9KEgWpajpeZMABvkgck0AYxBFc2cPxaPpIdmmretCxcWcVB9
MUsRJFsyf1X1YGBRAskWpRx4ohwHL1crOh2gjtLmyOO/6rGEM3HMzNBNC9ChZU5pxfZFQ3Ew6p1K
grkCm0RNf+zmZ0eFmbius8D36NYoTUK3444qhUaWSbDMNwOoZwYWC31VTEonDlrNggKY+j0/rzox
B/PwMavj3mSKINtb+Al7L8TdFr/slBaEU1+MR+a0iebinXKtoRoe6u2ulOM3eAqG7dOTz7+XQoOw
FlnEg87M5tdApwTPdgCAZsEHtpCT/FVgpnIbE5aMRg+ebQn7fa9/Zoh0tYwIT1btjEQnlUla0wEV
ynvtIkuuKGXhiGZIOuqTpCsM/rD/3S2b0ASO8VIDoVq1gq9pePvacscSQKrDoiM3SkQlQtZmc/mW
kyBolM373+4UtDqGI1Pz9Hz0gjOhCfuCd5PQ8zN+xVCmnawQT9f9CB5HFjMXmVsUWoocPYLU/2zV
6pMoIMQDr76+K5d7oS+LYjBm/QiEnMqXo50uP0O54GeIjzCuTkpXiRPZ5d3EobvKHkyUdYThyzs4
l1T/wcUL4Lx92jt+w0VDuomraRB46yhcPlUYIOKLzBLFM9ns5Xs7oI8jWsg+KD6o5Sc6vPZ6YM8+
mo5xUw0C2dmfKl/h7fRS8Ngj91jGPJJGFIxwgQ8KU9Ibuox7q4Q9LbDoeGvVAniPLlnHe+QzdkLM
BBafE4F+5YXlaF0WubFvZ8w87KrtUK7Wr+PbeCLxpof7ucQ+JH8gynqkuQNeWo37go08AbwDkYm2
j/iX6+EpUj4PQOPnsEbufxpPbw84ecV34xip6hiXi2T/CCjft4qQ6C2cLkXy4ovNORICLWN/Pgvj
F45n3nBxQ9cu8xrCkvgLuVXGblYvBO0noem5tNvYU419D3kdWPGzuC3EkEDUka7vKMeMiiZ/QHpt
qwhrDuCPhwTLB4qlNrN6qcJ1P0tN9wEfyVUdAm0r3raU9KC3++I8vDtwSOLLd2Z1xFFfjd7UBlge
QCUu7jmxAWO+iyMopvWuPOiGN/H3eQvIdJ6Ne6WYYW+xKlkEWzhTJXH+ek3pzr+cejQe0+6Mh93p
mRVLuoiSU6XOr7jU2zOKshF9CWgGjTc10Dd8QFSLYtNRCPB5NVac/uzZDzXA7n1bhwwYLaEgcEfr
QPk7yZQgrSU7H3RWiFPAI2W/a8DS9e5tfl0yq8tUxseBM6KKrP4R3ihZsS28sHbd7WGPjRAa7Ex2
klhd/zm4uKUtuuRud7K7Nui4MknZQmErXkElJyTgAMqGvXG/PiTrb0snOUaWgzaJJf9VHYI9Jvtj
30WOy6jhgmSs0blPDeGx/f/qjcIXqzSR6H5r/qduC7gYM5RntYmWPuz7EoqOj1gIMVs6cBeBn850
UCNa8TeMVlHd63iScZBTyKVVM5QTaruMGj2gnzWXanm/7H6Waoxy7cNUxNNF2ECRlzMVg73U5pWZ
7IpO9eqH0jLfNpDF0HixJIK5aWD0e+89hgQ64LQhZF5APcrIXydSvLVpiTsLb6fUfqgnJTb6ZvQd
eHQv/w/gDzoT/GaTC3LOcSL/jUGAKpBTR3kiV+dnmpMu1uEZPUtzWKSrqO/uyXVTf6YWUScCALLy
eoLjson4Atx1/4d/OTSPxhhFbGtkZ+FALQZ5s4NQUoDiih80/jbHQm5tQoxKYWN4lAxvG5z5F/q4
9xqbSCydHX9hXqu2uUe7JficOz79aiNc7JBrGNn37hZogAX53/rBn/ZbTmHKUi9Zw3ayPNwwBzrt
kRGf8+Qeg2wsLL0szYJrvnf1x98zllLsbpuA++HTbSW3VRBeA0hj+r6UzvS9qOUtNDPqUVfnWudc
rUTDsviqUcmZlkpbx1ggJRYLTwiA/calR3JKgZkfgiLcFRAQKJgRwYyQmVBwcibaZOtm2xOSsiUc
v3ZXU0ZZ9UKiWBfHi1j3K1XnNlZdG430+j0LLwKmIsSA/wUGzFxus3Oyy7oBwWrPWT15dF+bcRYn
Q0nsL9QuiYzMnontueoGcS2KSVOVi4AAjHOuUkwdWCQU32H49sZuAID2ol89pVCc5qREgmVj0zua
BKH6cYveAQH0U2W6v6FX6Qs2NTHuCAX5r5mWZ8H8+DlqJVFKEw5P/VapZj5YKP+t3QKkcrmrqtFz
rXOPPU2fWOe/fssh60NWfvWUuCoRjEulnXMMKO8G+1fE3OhZ/GeWNKTq2bJ2UFl6tBZgGhRuPLl1
9zQO3cv82G9lgvQjgxP18yjF7bgdYi+Jyw2h8mSuAuveJ1S7NqQUmX5c0pRy2ZAWpXBK3QLo9PBY
6W0tuJbtqLB8omLd3oSVBjkl3t02V/HR15y1kUa6u5Y4EMvO/U+vWPK8GbPfT9d13QZbB2tY4rs2
eaQ9gkk6NzVOTXstPfOR2rrczVJHGLideacUaiwbyD+xaAfKqjIMPXmvEHrz7YV1HCXZmij8+o0d
Tb5HrgoyLpOq1wUqvT56Sb7r7by0RU0SggJR7u+uByaHf6qORNdSaFBV3GjtR+PIyCiCifvirv0Z
9gCRDNVMHFKFixnV826Mmyc/AJY++Fea4tDe/DwRK7Up5BFP/oXEC2x2cjnZ1cs2FGvdzAYF4WtH
KRBZFtkW7G/Hjt29awSDT8iwpDF78issy88DiHm7Uq5xXLSqMXCRud00Grt3Y2v0AkRHt3V6K7zf
UQlaJR8ck+QRQ1K1rET3AHxMLD7FN+c09HmMm4KZdqc0RomCREe44eMgBwzjlnslzhhR/ETZya0i
koqFwYYpTluW05UDV3VbJVADsyRUGkjDgFlEriyoWuKtdnuIGihIPxkap6uVqrmgVPgq2860D8KM
gr7yGhaEzX9dBwfu64rK3537UXVq8f6XG9KU951ItfpcKoIWkIpHsyrNiiARj5nHS4uM06OmfYSa
XpJExPmYF8J4JyEWntlGK7u4sHvozwDttKe98d3ly0Cbmz4rQouVPaAjZfWC8I0/ds7q2hBtpYW1
8qo4GrAYpLtVTJ6iiGUuNMbRNwovXtQcDZi8sez/9l/IsMa7HtIbPYai6mC6eZTjKeDUFmcC0Xsq
83bSbHPWIPARCr8z3IZksE2Hkcta+E1WOr0s0WYE0Zln9kpbUkvekP22WxJfSPN1J1h6gEYumx4/
cJsaOjSX61QDYpbwnML6qbrj48pv/eDVRaHiQGWW9VT2FQJl3zRNOQtRZB9hA2ckQbv2QtKX6oZc
SAaupIvQx+UPgoY2+KDeu66E7VAtgu2ZdR8dllYM9KewfFjIAw2bjmV2sAonbPAKbcjGwoUrXNMv
+uvmcEE5uNi1hOHcAoYC7+g42rSgFFf0w9B2sxNAlrmox910bPBcDUIAUqWnexLfUn7ovFCJam8y
4OtErIc1jfD4ZH1eOap+cGPhtG6hCzAR+hQZ4QQav+Oh/J2j45pWs7ec4awVMFcGjTBhX9MhwyNf
xGh3oynE0Y78PGKL8N9I5R2BA06SFD/QWB1FKClJhdHGtTugBc0cWDRLidn2CTCk5TBP+xs8Otqx
yeXW8PiPyWbIBL+sOy3E5qf/9obNrxE1nxwN2LyBAScrCo6Alp8Q5hajhRees5UZjjc5I9azsxsP
ZeoX9bBCeoouxuvMPL2bemrkT/E3BX7wYxVomX7NhHdCQ/JTCeL7F2BHV8RgzAZHcscTf2fLupc6
om7SCPgRGNtB9YoRNXi9pzLMFDuuoszS7UW/PBxcHvJLKdmqxyrVVXYDDzcT4QlIIPy8N46zut0A
ioKgDRxqIXIbOjTZF5wMLy/7K+Tg1pIvHVx1hipULFfIZLDj/5Ass6FM3Y8n7RSpGUX22DVhc8AL
+LYLfyo3PIGk6gvfBOF3batBi+nadaTB6zZ3i+p4R9vGPi7XGWrdyY7SFbeZk3H62YOsEu8K4cFO
ogZ4k8ecRm73aV2QTawd7t8gdFCRg6bn9k2Rxzf02CsP0vD1LgCOaAgNRlDV2dqFVyOMHPLzGcRg
LBwKF1Ad/By6aIMYYUF7+bQnAGC2KlPmhYpbdj5O1Xx2xPz7/vXYY4QH2qofFTycV/YAl+OZ+cwa
JNrEPXyJKJ6CDIUaD7983mKnsGYecX0SLvKvGtCTF1r6lrJAxraL7wqHq6QYpaUrXRw/OsbReM+p
FXHc0jojtuXXUsI0T9jmcU7A5zjZyWmApB6IUU6vPMtXDLtBL1/XwCvwtEdMF2smleBiu0VUSd06
yMe7SytAShh+6NQ8QTr0B+4piVl5TjGijMIbI6MNUAFZ8ae9wjmgTM9LL/1ExhzCQWmlvIsRuoP7
MLhYQp5knOT/XfVCJnqIufXAXLPSqxAtS/tY1+E2BNi/Q5WPg7/0BPKDzLenQfg91JbRP08G9TfW
vECJq1g37ryALNQdNjyzHA2OYOBJSUR359W7n+HoIpfYgUbLcNx/LYt9RoxdluQ2/BccdXQFmf1Y
dUpMr57cXx462kxPGA4cq76pgmwEhambYOFTQmXNsRZnnB7IrYbIeyaeVx8p+G2yN1TJSM9jXuXt
bYITGJ6J/Xvj4AqweCwPwa78cMPV33QY8C9H4V7YP7z+/kIt5USOdQmjicgNKJ7vDzPmlMKnj0gK
U9VneW9UdPhjolsqUsLw+sd+jY3sks1gePPoC/SJ7Kigrkk/mn5EaqegF+x0DxgKUsfD7Yp3ot6e
gm8dgW6+IMRFebVP+GdHLpivtmgPxUgWLkCfw1Zo/T5818CV+nhTlvgfVzpHlNid3JQQeCCdErdG
xuLRCqwDO2jC4k1uvuCM1GqqEtVm1A1dY5Mu5M1VR0q2sZMux/HBdIPkr0wzOFMAI672BXyzBKfv
JBDM3NiNzW8PLs4ZZTNkXv7WOvlZUAkKBoY2Su9ORBpkTlrnONHJwMWR1byAvfgEMVBQgZwYh3Ou
WyoVGwmaw8Sx/Hy6hVa3gepYa+8FSglqCh9OWQQgwA1Wm09Zg9td6G45HS8yLq+1AH5SYCignnrt
OIhMURDTqXsyuxqZyT0G/qPs86gaH1eJtxyDYFA5/PnFhCQ29+/g7yOkhStS8YZVOS1kYn7GO9jC
j5n1JCjlI9yt2npcrJ3DwoWPkYlC+teN3DOXt9Wh6F5J/Urh2aRX8qf372t1fFPduj6q214HD5f9
Ru8pfVH8v7Dh9cHX+g10bsZic9giNfOUb0vQxAoR7zuqL0TZnLLnugIxaia5uaxkFHfZb9uk3/tw
ZZZAWBU5vnVgRPl4v7gcG+F10u7nuXBOENS1u3g+4rq8RtTXImzhHx2QQ55BT1u+kZ4ONy7HemWr
M2b+LmFPdEz2VDDk0uTiNJ4xZ1oaYx7XjGWek5USmUUGFfZZQ7er7t+q46rbmpljhq9Ztxu2kd5M
x8u2DrYyaZdRBA8VoKBWRwH6Ilm776YOFteLOUUzAyug3xUYlh8veKMY71pWanklr0ZiAOIbOmUh
QzURc4sQmHpPWQYmXxCXcmB+tMNKfp9rUjsCPMHzPrPjHMckXYAcMD8zPn6Hbaiw+dJ4MPWxuPNx
sKAUBgmIY96gPSxy/HMz9dnTfMqmhG1TOYlImNNo6/ebOGkne/KO8uGnNo6ha/II3EEmHe/26WBw
wX+S1RhtRpGBGJsUp4dPeU4brVO6mtUcqJ1kk7fZ3qgq8XKD52UuOatk6cVpKmXYxNR16r/3JYpQ
RISIo1bofmSqz9dcSDfHMBlZOYUiI/2j3NQCk4ubf8Nnk/TCWa5LSEmbCpr4vUcP8n9XPAsZMuz2
m8/eHb67IOchmB26y1QB7GBd8A8Y63Y5XDdKrtIs1hXjz3lI44GsXE7SEBNNC6MjuuKiVX845qg0
vzqM9r3BvnJ6/unLEYw/o+66sG15rNphpIMY7t9S/C5E2wXOKko9pnTyT5WRTTBRYd6xII6fc5jC
yLnn98lTR1MMoESnM5MtWr9BQoT6E4Lz0t8N+jhUTbLrFwRqFlPcLtX9ofbiJy4D4D+l/HF5dRmy
V+eIms8QHtGHxs1KkYnkRaG5JzhSLIyiZnXALphQPVMFQ3CpweUpJD5wniuvhv8G+PCWEukOvtmD
wkp/8hy5kqoyLQU4YVecD3VSHldd15ZcVxdwSYcVguwpOapAz2AZJVMJ/MDQuV4Q+ODnb7nY3kLZ
8Cjp+z5Eh2bTisZq61bNEZ/fR1BK/PGvdvk0VjdXwzE4B+iuPmSGttJ6T9DXn0uS5JK4Xgk+dfBc
TVM3RgeI6Sa+ZaOCNOO4Dga/gGaX5RqDUOY0VQTy/pQgDYuAkBPogrUHJNLQwj7i7JQbE2MXiWv+
CdToMYOUDUTt52ts1ss4oubjq/Z2ffDPLXghtZpA8PW31UkkwwVwcMFfh/UBmaboRymjyUCekQ3E
z/j+4/F9vnY7xrgwQ6tOLqfAW6qF+5vCVpJ4PT3ZCRXUjW5/Hw3P9lol4++bUcH2f+K3pIYd0Sdd
ZHEV2+lKWLPjD5MT9itHndFx2DxJMe8aumd7iv4xfuAlZsN473kRea8io9lOuw4n1nlAYPAKib5y
69bCeIXQGh+kRDnJuJ4FsXNWa/n+L7QuigQp2MlJrwZnxEe2wHVY1WF6CydbFVdlWmdn1coRsJTG
SHIRcipBMtY+kBdqnrE3D++nv+D4JU9M63YrGc0YX781weGabTD2GJYI6KbtiI4cBabmhqNVnMRP
KttVrA1/3aegUGiyJ+7HBKd444NjsJY0D1Uh1VqJPQKGOVRXbV2jnhIhGsRY585wgfFNduOjX1sY
4JNS8A8Y5KEQwXvFmjXQNiru/+NvyIaMImGmKkTd8Qzsm0Gb1Rpm229vI6ddPe0qVgoohOfTY3yP
7dZPBb3lrF8ewpHj7rx29CZcydMVwMtrQUZzkmuN58XSSkDz6XdfaLmicb1AwiKDNIUdoFBC4jy7
wwpxARn4HiYJ6mcy9cEfhP8WYqrgbFIwIBbwI1U1KNSpQRE/ZZsvNbqXxcd9uXaJQYEv9UwDDxOm
y8RnzM2hbD3i/WVikBW1v7CtEtuBLGXdOiQ/b9K7F/KFvQlstQb2FLZ+gnsXXC0hw8pSOFeTdP3K
Q8Px2CRwOXIrwMc6Nw4p3hgEVwyyoSUoEpt9zHRnmebhqtdZmkbBuo1IrCDgianOkr8Ll+WzD9ZH
FpPLskpKecOHXxmmi3nBPdQHheJb7h+XKvY/LhdNPfbpsmCoSYNZ3geXU2wdskAR+TyTwmQX0KMB
XQMHdAdnWgabpqMelYmvWQuDlXCDPx9Agg7nU8wlqUdXel36tk2ys9QjtdcnlVnCvRl+VuCyniWk
aa9kabBh4lIw0sA2Y8VGNsJNZlFWUiunfFfGTM09+BIexWM0Mf+RpLssbcKanVxrA4jRLJ38+F4z
lwACeCHRS61WlOlLRU66meIz41NBXHkJz0Cp1WOSAbkct7S9+oWTqaYzmZ3NNhMDj26ThmiRmOsi
fr6hdxwH+1oJBYEOJIQsu0sp74PiHHTHeMpW7R5kadH5PFMoF9OJh7vZ07bl/mMK+h+hcXUqLlY7
BsfAnY/hP3Au7nl3Ne3cTJG5IdghlS/92qUvrz/JpFqLOk9iYOlfgRw9xtzGTe+MTFMpf0P+pQD9
8HoAWamfgtJ6xrY/aonquYMay5TrZ0qyx66yr4aMy6oYVEBfcsXEcR/uIsp4xf29FOryqCm5ttCE
eOgkJHVHvrs+5kfWHkuvTCMnkWi4ZzvCfE6fnoVK/cYlxWRnMLRAnhLvODFG+hK94T1Oq03MkKdT
bY68VEMePnIme5MBfElkBY2MAV/9ZH5Bj/9ewHxIoNUYScuuZxIGV2WpmFhLsbDKI8xwkvCkMTU4
/0+LEVyNHmtBx0RNQjKoD1MYVgirOrlRD6Yx3toE0cAZYVL8ksCfwSBEbR5jNVKuymODc7IXoQRn
/nNS56r3xUxYP7DEFMn4+ds2tLU2AjpMASdBQfm22+Vcjz3bImC3cdAZox+Vx6Lv2oz9kcQ1XTK7
JsA8BI5eJi+ddL77FN8TeADJdKmmr7MEZUOXDPTZNNl9jdHJJJbvG8G2GygxE97WDnmvoc4gHC4l
kuKBHr3hKjMgbTujmeJ+bysfgoJXILu2Up1Ho4jWpo4tDK/FGImOmaOIPPmLJ1rDPFgXO8cZPQPk
t8xLs1sOjXHD8wwzXDAX7LoOxD47Oa9v1DirSoADGUvAuOrs/yQkPa0+H+IyWXifWohPLKYJ64rS
7c9axUaBv3pGG0IHXULH0beLV/XgCoTsD0KBC17+byu/ojkiVjXpt7Q4Y5tG/rDrtHr7Jvh7KrJJ
IhS3o8reXvMKyge0ocaDJmf+73p/EGb3SVKSaXgfVi7CyOOzQmbHDFESmvF3l4fzxv8SHLhyniAi
UaaM/U+JZvaGcavRi0Yb6riDKr3maRrgN04OsDn7w8bXUM+oEEKflEgkb5yuTOE9Y48LibdOzhP/
eVswhl7UHp1zrL59SIlOWvoOeaidpad96CGhfvchN37xX1rP3MTzVOyEREZMhpC1EdyQMbs8D2iz
2w7BYGKGLvGJHGxz7n8kPgNRTsUp56ZAH7JUZktoMCHFPjRsk9rmXM1OFrJc/CQSc/X0HDWoFQGJ
kr4Pt+wU5+3uvjkpBz5aRyu8idgp7ypyrY2d7QbAj9x5e5x5rxiuXKd33SpZTIXVCOrMO1Ms4qd4
wcHKgs0zOKmk1BFwnLDs8diw7j4vav53D3ex0rPwVn4mTT7tmiY/Fjp4WnM+Bxmc4NxGQBfK928v
MeCXaGMVu9lqoLNY8Igae7wpwEoYMbeLkeh8Y+x5wx9zH8fshZVjxLRh3BDrqHpUBS6Eo7J/SCFZ
KIN68OrK+3gxDWTBfWCE2e+hIow0NXAJ/1bHqznyOjgfeUyUqyEE++NqAiyky6U8Xj+qsj0sVuuE
O/Xf4OS9ynnQVPtCZlTEDlS5WTYfnXbhzDm6vQQinkuv0JDD2kLCG9N1MnecWdiRgm3tQ2onvlOa
SFoa1hHgZMRXfiknnVpG2bUCfNr98zqDJV5VJXgzDXjzwePDShtRhF1oCcFRyup1O/PxRtUdpD1y
5QfPMHggyU6nteD2bH8s6+BbyvxpoioSCQevT81eF7yG6veXyyPvm85XSo7rbvh4opJzfiXV9yhb
FmCiodKlIWyLT+/y2XU6/wPaCBsZqeT+0G+JdkwvZspoH8qp44K5IXJ3ts+PczegjMO5Txqq+2MH
igyE4kJZoPYMFKbUJjGYTO140jBKXpPAMgxjj/woiko1ozwCBj+jgsgt9GLOvwaqyG5PiwjY80cg
WRcQwfgP/TfiuszRpxY9ctdKnSLu7Yfhy8knEW6UyiXjiBcMINtlJVT2nIo0WUMke88To7FBe+lg
5g9SuqCo7c1d+Ssp4mvWAYQt3CY1E6tNnKJ2VwKFcLr23TjqZMIkcuZL3VVeoQmx4Y8oG1T1lBRZ
/fN8S9Btn3I6ny+m1eyNjMZlOkgWh4JxwwD+AwXPlKnEFnTdjxKGNwAjjWbOkS54ci6XFCDtRf4w
aZn4rVR/YhJZ+5YQBWCHn3++5aSgws2grwotYKXql7WiTKIy1y0RPoWpMaEo7fRdQ6knqUASJbtZ
yRDET6X5LnJgo18hckIoN7YYGoIQdhPnhD+li80YWI/MVN7DcTmoiK2VvtCwYjub+ppOOpURUi1Z
uS47apJz/LfV6i84AImQ9hIiLLFvZCd7Y/lxvlU+jHHZgj4oYhR46yMoqptFK8FdqDx3ZwmrJZVb
BE0achRyjWLu3Qr718Lwn0vFnIMhJvbmvJn1FB3irD9Ad3xfWXyT0hzUmy/tGX8EbCfJ6M8iGvCC
B/mTxtdkHMghZPOJqW2RFXZfQaLiPYwZV6vQviHGy1NvmkWX2lN4QI6rMJ7moBPrz0q1Gby0Kqi9
NTQikCq8NdgoITYHKaUURoRt0XjzTAbnsB2K236/GyhspTlsMJOlX3D9UIDnD776NwBkqjleVqaA
88EkQDZs/9wyEEICx0wnT+degUBGKy/6TxfdnQoNQChWpL2qHNvaGTsJ1UFYHlWpXk7gDEx3Yunu
LBcldv5Is4bbeJstolMATzBwxmMcyvJeCijJAX/gPCGt3LZK2nCTYidmyWNO8UjOjKfCaAWEloD1
rM85Sw9x2283cy+M2uaATFv+Ils8o3kgc+ry7r12PORi3k3nzD5XnBiq7Hz6qY/pqTBVMvpck3+z
MrkN++d25+9q2EQl/h6ubL/vODam7TgQUfCzTHPNMB7Q+rIP8hw2B9gXf5NajDSkp8IATtiiaOo3
TNFNhWqXnuKKixXSnMQD+zW+IfqF280ndXSTRyFEX5+Li62gZvtYdsb/6o3bl3pWiqRqCV2V1Vxb
2S2iKzC8nhXIil67AaWnc+sEXTZqmYsbnIwaH9YVEWT/kWcV2mv+oIrlzLg+zX3Q3SIistcCgKR/
8CjIIrHTk3X6hYUV7Pe7X3hvdX8eJy0x47bTq44Bv61w31HLeMoj0hcJV2vitT0hbgH6qY3FiALY
FfF/AL4NHyTlCzw9iklfkub2/SknBV6i27yNey3xnA6OfUE1QwT/bnDQfZAS/4KLCGsVcavpb4El
bWrT0zC8iZdUXQMRj1pOFd/j9TSEL/0Mzec/52LnTofuw96FCilMvKROusYTP7/vRIxJjZwp9pA2
ze5mGjw4J8P5+GWvAlG/9esgpWOBXqyelC5NOYaPLLsnvUS79Ps8abU7CIDCgsUayyJBSbhfgw5X
3IeO+vYf3q7bU4QqCHDeOkiv5Vzg0kM4GUDgAluhLC318BIahpnNNeOsbP34W/DSwZjqcztz5N3j
VbxyUD4CM412fNO+U4HhtkXcMuSF5iHke2zJErSQXYnEX5+lg3WoaOJdlGNmyab+wWZDO++PMKk2
nBDsEVlwXmZ3/gfy+4JmthGget8cD+KdxRUcp6SpX+3ZEO3DeCzBmnijuy4muD7i0V/NzmA33hn2
4vEqT6Iw/QaheV4xMk12oaVtN7gCskeey9DJiibRsPArtxIm6/M5/CComRhHt9hvgNDtGw8P2FMr
gHuXiJbLKQpI1EZ3ziKXlQS2jKGzYdKhOJ3S+s68mF+nCvW5H7S9Ru2URuVjyb3RRgWexLsQcA9h
NCK5paeNEFS+DWdkC7w58aE2QaRGvr8W6NEnXpqYRMqvoy6KR9UPq62PCeIm96THzgoNxRTMPFl/
sjuZE6xs03RDDStAS39fyKw2e71dGPVVwGdU4PcUI8avcqXrCQOvG1cbkBSXcVSUySkW9lTXy8Uv
ygvg8tzyuBbcyDq5rSXjPv9yIjnxSSdaO/jVl+rvMhj11GLxUvlMwZQoE1awxQ1Lg6sey0ib9c4p
UCgL5Idq/LQ5KxcfyfV0RGKg7dsO9dJEj54ASKlK17/JvBWJ0icLFcUuvx39PN8NOQc+AaPdBkgJ
0f5UnpIAZo0gUaRg/ygWNVChp2oWlnr1b4ZYvpSBVZuhVejU1/OAlozoHXSC2/Ne4DeS857xbIYV
8CUe/BMfzcbbW6G/2WSPsh18IHnoNJrBQj66mRuwPzRE0Q5X9pxVqkktBZaWyWO5KDENvKeqPkYP
e7jY10lUao+9dzl613xBImCTVq7ES3L6u/GQx9o9DbtsfPMFm2GDVAfq9OzY3KC/1RBfsGjwEe9s
H2Yt7jD3DQwzV2VcM8xwsJlpCUfDZfyY1dLUfUH1ki3S48UODWAu2GoENvsYQImDdBcrmJ9TsWPC
kpjsnxPI46H9PWks+PQIfh2lcxaVtkuRA16GRdMF6bZEGNoFErtQkM/SrSmd2Pggg0CLdZcjGr79
AQpV4iNrG4X52qxoElFYpYrKnuINq9YeInRs/IstRUaal7l9f6nFVqQ4M9httl65lKPTlzeZgYzW
jzfnjYPuSW35xCHJYgTM0bvIJJTOpdbvWVfkNsbnoS51MaVDhb499pQAyHO7Wp7EoSLefmRutigS
7K1UQz+Kco+CRiZlUnma93vqScq8Ex4ar1Xa1iziv6mwMLmklpJWg1UJTZzAqGTmT73+IMyfGkZW
rkkub4GrHrCMXyv+wgaROx3knWZEFQU+9ENnhm8KjsTdnotvxiRv4fJue0TvF2Lwc1pfPfBLBe1T
f4IspF0qY0/SrjBFbnmTsztu+vDPxZ3vH+lt2dMXmaQhfN8SlNZnPkfSh2YPCMaOZz8LiS2+oP+R
mMsmfP4r3Fc8Qk9tYbsNzEnFakc0Tqv6aZebixf2HBltFVnZzceOD6RTdsPWJWM6A1hGEJaS7qkG
eJOyybpPGVKaJizPW+5+3ZPl4wetKahlpUmiddX8dVrp4TH8NxL/bJ5i0TAiVJF5iLP219HyWeFK
mtOoOCg9MrAt55CjPTK/TC7Bzx0W0Y72AzHcVGwKPDkqgIT4nYCzEJWy+6hthVhNumXRdHzKMM9e
A2yiieR5opTPEGsA5rSeF5Vf7zNMuPkLs6UiRmGkhejxfALypb5QBV8lZr6nZKvlrT/Glc+DCITn
nVS47+pnKH9xD3QHrIh0HjbaFd8yqT5nMmuE2jiFd8Fr47IJT+EVNNwE17oqIU8K1RzM8M6kIF6w
nxfWwe0AjueSHh8l7iBrcp9YVS0z67rNemohHb1Xju80ySDJSua0nzrHJIA0utSEO6PTyScVsD0c
aUmDe4HPNLjqU/nkdKcJ498ATBwkWsJ67Nf+G7N1Luutw48Kkd4zp1zhQALBWl0f7HIgUiHGmerC
k4dQBy2jhawR2vBRDax2h8QSAehU730dZB+p4ZNFYztW9wotlHTBFk5UwFCX59MHz3J0xgELPNVi
0wXrzMfOCxlLF3WubEFAGHDqeoIuyQnq8uObZk+LGK7skupYLY/heLaAFOwO3NYklWapETWwc/Gk
ZL9/TweCBiv65hmTQCq3b+inc2O+wqB4Jxq4Rbvph7ss/sEfBM41WRkAg8CABtQo2gS8K0OgAilw
/GFMVCnJmP8993LKUcwjEo09j2L8NKiuc5qEiycI9mZWX9vaBSxZ+Y2t0Y8GXRFZ/Jj1Lgq15VJb
GWDPw00TkhP5l26cnzqWMvEmecpM0oi6bOmx19O1lrzojMqO4vQSBX+0gQAFbWRc4QvuIxQJLpSD
B/X1t5K59+Lwz1hhoWIQxX2f5aK1EgjcBViSO8iGXEoT9UxW2TqP5/0YZxEJ7IKbabtsLopqTC8O
YcgMS9pFZSzEl8WCPhjY3QCnEN4eDkaadCLeeW1oHHL+dI/FTKdzYGhGGfn+XDM3LtEXto7wIacU
HRHIobeXagCZ47LD7rvMvLe0PhFcoJrRJXAQHRDUoyo/+J9F8rd7AnYWbn+yy0Mbsxq2Q3wB9eCu
BEI/hHwcP3n1o5DE7BWvBuuaP2VoNR0qa7t/xH8hmO6izIEVHfmdfmeCWsSZlqdBdujPk+7lDsPy
UTmbEaiA2SpYaTpUvIZn5Rv5pHmpXzOMfDB3A6y3QUf5MV/oXPCnslc1yD3ZfTo9e/VUTlEfyq7K
T5n9NBmXGegZo9veSI/4ZT0Zg8Z0kp4bcQWxLi+EP0KtiETLw+Rh4Ok/n9AvuCNwWz5JncOyF0nb
KbwqD/8HsC5m1+BlByQfpdo9Y1udwoYT5IGZpSd3Owe+BTJYGQZoarhbpoVAyt5W+DxX2+dw4lfN
K9wsmXeDGz+fUXvT2+La1PkrGha/f1cskma3LbzrOCzwU+aHfRiloQngarBslHGy/WOLkN9poARQ
ZgrFZ0xrHeM2w2h5qw5be9dkvLxA7sDfvQbHDKKRjKiPDa145kum6zRt06kNf0EfDs9HV9vt0JBf
kFJQRuiCWZKlip94ALx4l9YV8s5LlPc1vr5N7HeYykfW+dYEEbhatuzUCDYMcuS2ZBaqadORvwAV
v3zZITnLiEYUwjdbgCCPj1phNfzr7+pWL5X3Oaqcsy8uYhi3GyGEivhyFlC00jabriRnKW4ASb+u
PAti50DNI6nr8UNXbKWz20JXvdpKDaufqhlXSQou406G0P6KBYLm
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw5a;
use gw5a.components.all;

entity UART_MASTER_Top is
port(
  I_CLK :  in std_logic;
  I_RESETN :  in std_logic;
  I_TX_EN :  in std_logic;
  I_WADDR :  in std_logic_vector(2 downto 0);
  I_WDATA :  in std_logic_vector(7 downto 0);
  I_RX_EN :  in std_logic;
  I_RADDR :  in std_logic_vector(2 downto 0);
  O_RDATA :  out std_logic_vector(7 downto 0);
  SIN :  in std_logic;
  RxRDYn :  out std_logic;
  SOUT :  out std_logic;
  TxRDYn :  out std_logic;
  DDIS :  out std_logic;
  INTR :  out std_logic;
  DCDn :  in std_logic;
  CTSn :  in std_logic;
  DSRn :  in std_logic;
  RIn :  in std_logic;
  DTRn :  out std_logic;
  RTSn :  out std_logic);
end UART_MASTER_Top;
architecture beh of UART_MASTER_Top is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
component \~uart_master.UART_MASTER_Top\
port(
  I_CLK: in std_logic;
  I_RX_EN: in std_logic;
  VCC_0: in std_logic;
  I_TX_EN: in std_logic;
  I_RESETN: in std_logic;
  DSRn: in std_logic;
  DCDn: in std_logic;
  RIn: in std_logic;
  CTSn: in std_logic;
  SIN: in std_logic;
  GND_0: in std_logic;
  I_WDATA : in std_logic_vector(7 downto 0);
  I_WADDR : in std_logic_vector(2 downto 0);
  I_RADDR : in std_logic_vector(2 downto 0);
  TxRDYn: out std_logic;
  RxRDYn: out std_logic;
  INTR: out std_logic;
  DDIS: out std_logic;
  DTRn: out std_logic;
  RTSn: out std_logic;
  SOUT: out std_logic;
  O_RDATA : out std_logic_vector(7 downto 0));
end component;
begin
GND_s14: GND
port map (
  G => GND_0);
VCC_s5: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
i4: \~uart_master.UART_MASTER_Top\
port map(
  I_CLK => I_CLK,
  I_RX_EN => I_RX_EN,
  VCC_0 => VCC_0,
  I_TX_EN => I_TX_EN,
  I_RESETN => I_RESETN,
  DSRn => DSRn,
  DCDn => DCDn,
  RIn => RIn,
  CTSn => CTSn,
  SIN => SIN,
  GND_0 => GND_0,
  I_WDATA(7 downto 0) => I_WDATA(7 downto 0),
  I_WADDR(2 downto 0) => I_WADDR(2 downto 0),
  I_RADDR(2 downto 0) => I_RADDR(2 downto 0),
  TxRDYn => TxRDYn,
  RxRDYn => RxRDYn,
  INTR => NN,
  DDIS => DDIS,
  DTRn => DTRn,
  RTSn => RTSn,
  SOUT => SOUT,
  O_RDATA(7 downto 0) => O_RDATA(7 downto 0));
  INTR <= NN;
end beh;
